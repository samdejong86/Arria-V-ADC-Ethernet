��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��N ˉjU���&�O�r�p�W�M� JK~��Ixh�5�����0�z3���`4�o���y�ȋ��:� �X�ct�'�.nj�����fPߴ`n�Dj"�}��?E�Y�q�U�H����#��\�}r)��K2�.i$Ϲɹ�$d���hZ��S���~��L�]�y<�7�����I������d��|h>W�nqC�?Ը[�v��zLχi)��y>#^�������&����#`��ۓ�Yx���	�� �4����nQr��#sUt$ �S�?�-�}V��2W�mY?��{a�
��Ŗ7Pn'��W�B��*9u�W
:�u��}���5��萊��f����m]K�@Z�����.�>�p��w�	K���`A�s�$Ӌ�CT��o|���n��p� ��0��KԽ?!�xn4�f�L�r��L�9�b6�t�����h���s7� �˘�ʇ����PȆ�
�^����ᒽ{���Gr�p����~�����h����x�2�ܴL�ܱ ��X0�
�n��C�i.x·�)�IH�e��7˺B�;[�ȋf�z4��?��N�r��)�^)
� ��Ț8�7!�D�/�0u&}�{�ŋ`��F��Xt"C<���	�	�7=.������!M�mM>I�f���8���є�ϑ어�0�B�jO#���#4%��&ĉd2�_H
�Ӏ�Z�e��@w1�J8�A���n��3<;�b'%����x���6w'����B3�yY��A��4�@Y`�?O�HVi��z,�E�?
��������dj�#&!N�z��)�4�I�cb��S��z$�#����Sů2��i��k`��/�?����̪Թb{'���xJ��-s��g<@�tѤD��˘�85޺��l�8�����^�˪�̿��(��=)���=v=}�z3�:�Ϊ0^��=s�Y|�=2B���}kJ�̻�\a���ɻ4^���o�p�*��\o;lQ<�� �������	��|�^�rK#ͽ�|�ܛ��KpI��D26���M��!�?�9�=����4=5~������n�6�Z�!��}��jo��#�0j�3R:��_�43����L���	��@y�(������dqs��(�=U_�e�>1�3ڕ\�؛�򧴂���-m��5�I_boh۶L����`
�5��	����ٕ�9��0	�B'i0GyB�	���F����a2^������<������F_u4ģ�+�n�R��Ǘ���6�o��8�r=�:�$G�
}k/�Q�sk�L�S���o�y��!���-��c�����X�h_��:��wɬ7���;�*v�6�.q}4��!j�?��:���L�Y���}'T���"��ZK�ȟ�r^���D#���D�C��D�=�x��s~������:��*.¡(�k{[4O�H؅��Ͼ�P72+��Jv�~����8J�� �Z'�����h������af�>��U�*c+9O���ܹrREDX���m�,����6aܙ%G����R@���-�L�}w[챿�p=w�x�����<Rۧx���+�r%}�ɍ�?�i1���*�����P�=(�9�������L,�@�8"�`�"w�p.�$n�j�����%�u�|<�dY������;�)�i���_�����u8�(�cI�#�.�ڡ�`�[���{�l~&���v�#"��]��5--�g�� �Y%���S!C1y!t��6�Z�D�>H��I��1kS��D�oST��EϹ��x)��Ŷ���_Q�!lD��߽����l�4���[�X+M[��9�g��`�b���^ֹefT��D�[����M�X6��,��{#���u��\���)�D�!����񰸝��3?����tS��s�l��}��Ԛ��[������ \�Ǐ�:g������mL��I�Ր7CoAf75�2�u7*�l��ߓj/�U�q6�	d�h�Mu��91p�o-��:Qu���l��k�=Ra�&�<�Zqc'+E��${�$��sP���e�uʐ�(F�Ĕϓ��r�u�4h��>q��Q\�-ӣڇ���[W�٬#�'�� ^�D� �RO�|�N��:m.D�X�@���xk�`�0�~X�F;����4�V2GW���A@X��Nov��A}V'�q\hU78{�BoI�pIH��Ä����������2��=�����Q���""&��q�6�3��<(-bj/�ϔ��S|����4
��ԏ�]�2Ѷ�\8�����{"�'6Fk���8�O�-0H g�9��ޮ�W4�V�1ߎ�yë� 4u=�}���$R��,F �ڦ��8�p��D�c��\�O�	�&�g�a�Ew�ȧ�����خ���$d�w�����@�)��Z{o5�nd{�P�	w�D~���~_�t�t�^�SF�$A��6���+m��s�/D�씲%��s}Qȇ/O����Zb��1��mH������v���<�~�>�:J�,�2�2 �s�IX/�p7g��i��(@� y�Ӕ��ETC�ϒ9�W`�^:q����E�2!��ג��iͩ�J�����߆�/�`>��`��)c���{20�$�-��������R�@cM��s������a.�T#�8�U�G�.�������5b��@������3�B}l�B��J�����i�-v��r���jJ���8�3��oE�u����b��g̕6���ۿp��T�t�j��׈�9�����L ���H����T�".$=Pǡ��I#�e�µ�{&��V ���u�d�_(�y�KP--s�'�/���3A<jB�	鋳���1m�^�$e6��Ӕ�2�8�3FPa��":�R�d5z�:�R�J7�l8m"��/H�Ք_��;��ȟ�J(I�[��U:�h�F� ��⬀��4��?U�;�n�����9x�a��.óeԜ��5��j���9r�s��aR�L��$�.Zy�|�-j]�T�óS6����*#��}�gzEl�~���t�-�t���?e�Lw�������IC.�r�����f����b,��4�>X�5�5׬���Imak������dL	Ǫ��:i�ֱ��
��OX��y�H�H�-ג7�Z@e���2�\���pN��y��N�,zweim.�Vs6�(q<���C�F8�>���㹯H��9:gb�u��q��Z8I9���#xI��KU�'͗��g��r�}�|��� m��d����y~
��ds�\��M0%J@�v�L|q�r�-ث�(A5d��6���V� ��#�ף�7t%�LwtRV����R�#��T���A{ȃ�p��1x��N~�����KTYbl�ҭ�-VTH��ރ�=�E�Y>��*7���{Sr���P+�Hv�Jo(T���-KL"b7`X�m��6�{+KzF���R��F�d�Я�.e��Lr������a6��.�:�Q�ry�	�v3���5�a����$*��wT�K�1�M���"�־)C��ʈ�p6(I�\<�Xy�C����\���]��f�魻�@]�u;�h�Te�����N*3�F���4�7��0��r���M���a$��w;�W,�!�Ӥ{��Z�9tSaȜ�J�W��3r=Q���j�GM@��fp�F��*���7��K��ˬ�����;3�����i���k��+q���Y���g6�{��+�紁]ʴ�æ��n\����	�gE�M׹�tΕ,�]�"��;��b��*���6�xl�?��3/�z?���	��'���[�I�+C�ip;�i[��$�4}��C��f�f���y#|��7�| ~���bw��D�����s3t���1i�Q5n��Aa�k;�pW��Y�͕���Sâؿ޻��Q�'�L��aNg}�&�'���Ŏ��X�B���]@�����z:�|x����c�͖�w똊r@x
��-�ۻb�F����D�r�l���1	;3p�"���ۆ�B�"�jl�M�Q��@�N��������>:B[;�ܖ�	��x,����P>6���aF���j��'s��|�@O.�F��
�mvSGf�@Z��	����D�(R�������^�+���|р$!{�	�%.�D���3�C��"�B��G>a�yrڋ+�1??���~˿"Cʅ�7?.0����tz�]���]%(#�<N��^�a`�Bd���>w�O1e�ip$Ԏ����i���425����fl�|L��7���֧�ZV�P����GH�)���#B1�5�T���q���_!�I3A�/�� /*kNj9����1�S�Wk��zsϢq�}6�zt(���W�@�?q�}-����>!�`�1�#���~2�'k��W1â�4�\�iB��G<K���5�}��C�y�������S�ۘ��c"�C�c�h:�&�B��� R(œo9,�f�!��Z����xج� V<�P#���i��'/Z5�I_�#�����o=�d�#�kg��s�PP��\��@��{ٺ��+�D���8�.��3�(�c�fox��h�3L��u�ػ{��mi�@%r�c�I�W�����k���Ж�D ��2���o�6g��q���2���Hc�>�� }/�d6���,�j;����H��ٱ �3�Àl��%��Z�λ�QJ�D�?��M"��T�K�^G�<����?��