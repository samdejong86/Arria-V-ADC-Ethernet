library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--my custom modules
library work;
use work.my_types_pkg.all;

entity ADC_testbench is
end ADC_testbench;

architecture behave of ADC_testbench is
	signal adcControl	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	signal a2da_data	: unsigned (13 DOWNTO 0);
	signal a2db_data	: unsigned (13 DOWNTO 0);
	signal CLOCK		: std_logic :='0';
	signal SampleNum	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	signal waveSample	: unsigned (15 DOWNTO 0);

	begin

	ADC_handle : entity work.ADC_handler PORT MAP (
		adcControl=>adcControl,
		a2da_data=>a2da_data,
		a2db_data=>a2db_data,
		sys_clk=>CLOCK,
		SampleNum=>SampleNum,
		waveSample=>waveSample
	);
	CLOCK <= not CLOCK after 10 ns;

	process is
		begin
		
			
			a2db_data<=to_unsigned(8054, a2db_data'length);
			a2da_data<=to_unsigned(0, a2da_data'length);
			adcControl<="00001110";
			SampleNum<="0000001111101001";
	
		wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8073, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8078, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8079, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11054, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13843, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11721, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9367, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8148, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7690, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7545, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7456, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7443, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7439, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7477, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7495, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7518, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7561, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7591, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7636, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7655, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7652, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7700, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7711, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7727, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7749, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7770, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7799, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7780, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7812, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7828, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7841, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7848, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7872, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7887, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7894, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7916, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7919, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7931, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7945, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7959, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7948, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8003, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7998, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8020, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8037, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8076, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11004, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13837, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11735, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9374, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8150, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7696, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7544, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7464, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7439, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7438, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7464, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7502, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7523, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7567, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7596, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7618, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7652, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7662, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7692, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7702, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7742, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7741, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7787, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7788, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7803, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7834, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7835, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7844, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7844, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7867, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7885, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7895, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7901, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7924, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7926, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7944, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7962, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7951, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7982, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8078, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10974, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13831, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11733, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9370, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8157, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7699, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7531, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7472, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7440, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7463, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7471, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7496, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7539, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7547, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7573, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7619, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7648, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7679, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7686, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7722, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7735, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7745, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7787, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7785, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7797, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7818, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7827, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7832, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7864, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7866, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7875, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7899, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7897, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7917, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7934, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7957, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7961, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7980, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7984, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7992, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8016, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8023, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8039, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8034, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8030, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8080, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8079, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10954, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13841, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11766, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9394, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8154, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7696, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7547, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7448, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7427, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7446, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7470, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7504, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7526, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7567, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7596, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7606, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7655, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7665, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7702, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7722, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7730, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7752, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7782, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7777, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7807, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7808, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7839, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7833, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7857, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7862, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7866, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7895, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7909, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7923, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7930, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7942, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7954, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7974, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7979, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7998, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7987, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8016, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8035, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8071, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10900, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13824, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11793, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9403, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8164, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7694, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7544, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7474, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7429, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7436, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7493, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7509, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7540, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7549, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7585, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7613, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7648, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7665, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7695, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7713, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7730, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7746, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7769, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7781, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7812, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7814, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7824, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7840, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7847, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7875, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7876, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7887, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7897, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7909, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7946, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7946, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7965, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7965, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7988, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7997, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8023, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8039, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10866, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13833, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11811, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9422, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8163, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7704, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7548, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7476, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7438, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7452, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7490, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7518, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7534, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7559, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7587, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7631, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7641, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7668, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7685, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7695, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7721, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7760, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7752, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7784, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7816, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7832, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7822, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7843, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7858, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7864, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7876, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7887, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7909, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7907, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7932, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7950, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7949, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7962, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7992, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8007, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8002, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8017, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8037, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10842, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13839, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11810, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9420, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8179, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7711, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7550, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7460, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7438, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7453, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7459, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7486, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7522, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7552, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7570, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7596, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7634, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7672, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7682, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7702, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7727, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7737, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7773, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7796, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7781, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7818, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7830, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7857, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7854, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7865, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7884, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7888, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7898, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7920, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7925, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7945, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7968, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7956, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7999, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8018, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8024, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8032, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8071, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8038, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10796, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13835, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11838, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9432, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8167, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7708, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7541, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7469, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7442, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7449, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7475, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7508, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7528, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7559, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7575, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7611, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7631, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7654, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7691, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7716, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7722, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7751, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7779, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7791, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7798, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7819, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7829, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7836, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7856, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7872, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7883, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7898, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7903, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7924, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7927, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7950, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7952, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7965, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7973, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8000, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8007, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8034, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8032, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8071, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8076, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8039, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10760, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13837, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11863, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9455, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8172, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7704, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7552, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7476, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7452, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7432, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7484, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7490, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7527, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7564, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7582, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7612, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7636, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7664, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7676, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7710, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7724, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7738, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7763, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7775, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7798, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7821, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7839, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7845, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7857, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7872, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7865, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7884, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7914, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7907, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7926, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7942, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7956, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7967, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7966, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8002, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8004, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8024, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8038, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8035, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8074, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10749, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13840, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11870, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9461, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8175, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7694, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7548, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7482, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7442, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7434, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7490, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7514, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7526, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7556, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7583, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7618, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7652, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7666, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7688, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7709, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7734, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7755, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7764, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7794, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7815, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7808, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7850, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7855, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7859, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7873, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7878, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7900, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7904, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7921, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7929, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7941, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7961, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7967, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7969, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7986, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8003, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8016, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8037, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10697, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13848, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11887, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9467, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8202, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7711, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7562, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7452, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7431, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7444, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7494, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7508, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7553, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7547, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7594, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7612, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7635, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7676, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7684, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7704, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7743, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7740, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7770, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7779, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7803, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7812, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7836, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7840, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7842, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7855, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7876, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7882, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7901, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7927, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7936, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7924, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7965, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7966, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7985, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7995, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8015, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8039, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8074, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10670, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13843, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11905, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9483, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8197, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7722, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7549, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7470, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7439, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7468, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7467, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7503, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7528, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7555, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7580, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7614, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7636, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7656, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7681, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7705, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7735, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7759, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7768, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7779, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7802, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7823, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7825, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7840, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7864, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7880, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7884, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7882, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7905, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7922, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7921, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7952, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7966, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7970, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7980, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7998, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8031, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8038, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8071, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8077, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10637, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13840, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11931, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9495, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8200, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7732, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7544, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7464, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7442, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7446, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7470, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7500, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7526, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7554, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7586, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7628, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7653, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7659, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7687, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7712, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8073, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8078, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8079, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11054, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13843, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11721, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9367, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8148, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7690, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7545, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7456, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7443, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7439, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7477, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7495, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7518, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7561, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7591, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7636, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7655, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7652, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7700, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7711, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7727, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7749, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7770, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7799, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7780, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7812, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7828, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7841, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7848, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7872, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7887, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7894, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7916, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7919, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7931, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7945, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7959, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7948, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8003, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7998, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8020, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8037, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8076, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11004, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13837, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11735, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9374, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8150, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7696, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7544, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7464, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7439, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7438, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7464, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7502, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7523, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7567, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7596, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7618, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7652, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7662, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7692, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7702, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7742, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7741, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7787, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7788, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7803, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7834, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7835, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7844, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7844, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7867, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7885, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7895, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7901, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7924, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7926, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7944, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7962, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7951, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7982, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8078, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10974, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13831, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11733, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9370, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8157, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7699, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7531, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7472, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7440, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7463, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7471, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7496, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7539, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7547, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7573, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7619, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7648, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7679, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7686, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7722, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7735, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7745, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7787, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7785, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7797, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7818, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7827, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7832, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7864, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7866, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7875, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7899, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7897, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7917, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7934, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7957, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7961, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7980, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7984, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7992, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8016, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8023, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8039, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8034, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8030, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8080, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8079, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10954, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13841, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11766, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9394, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8154, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7696, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7547, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7448, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7427, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7446, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7470, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7504, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7526, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7567, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7596, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7606, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7655, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7665, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7702, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7722, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7730, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7752, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7782, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7777, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7807, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7808, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7839, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7833, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7857, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7862, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7866, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7895, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7909, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7923, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7930, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7942, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7954, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7974, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7979, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7998, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7987, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8016, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8035, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8071, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10900, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13824, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11793, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9403, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8164, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7694, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7544, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7474, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7429, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7436, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7493, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7509, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7540, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7549, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7585, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7613, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7648, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7665, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7695, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7713, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7730, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7746, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7769, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7781, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7812, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7814, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7824, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7840, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7847, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7875, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7876, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7887, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7897, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7909, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7946, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7946, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7965, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7965, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7988, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7997, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8023, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8039, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10866, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13833, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11811, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9422, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8163, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7704, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7548, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7476, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7438, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7452, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7490, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7518, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7534, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7559, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7587, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7631, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7641, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7668, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7685, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7695, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7721, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7760, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7752, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7784, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7816, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7832, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7822, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7843, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7858, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7864, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7876, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7887, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7909, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7907, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7932, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7950, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7949, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7962, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7992, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8007, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8002, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8017, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8037, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10842, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13839, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11810, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9420, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8179, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7711, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7550, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7460, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7438, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7453, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7459, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7486, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7522, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7552, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7570, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7596, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7634, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7672, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7682, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7702, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7727, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7737, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7773, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7796, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7781, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7818, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7830, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7857, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7854, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7865, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7884, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7888, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7898, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7920, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7925, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7945, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7968, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7956, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7999, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8018, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8024, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8032, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8071, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8038, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10796, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13835, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11838, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9432, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8167, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7708, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7541, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7469, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7442, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7449, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7475, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7508, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7528, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7559, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7575, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7611, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7631, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7654, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7691, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7716, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7722, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7751, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7779, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7791, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7798, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7819, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7829, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7836, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7856, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7872, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7883, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7898, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7903, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7924, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7927, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7950, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7952, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7965, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7973, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8000, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8007, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8034, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8032, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8071, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8076, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8039, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10760, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13837, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11863, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9455, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8172, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7704, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7552, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7476, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7452, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7432, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7484, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7490, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7527, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7564, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7582, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7612, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7636, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7664, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7676, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7710, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7724, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7738, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7763, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7775, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7798, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7821, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7839, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7845, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7857, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7872, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7865, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7884, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7914, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7907, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7926, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7942, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7956, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7967, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7966, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8002, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8004, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8024, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8038, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8035, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8074, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10749, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13840, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11870, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9461, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8175, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7694, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7548, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7482, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7442, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7434, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7490, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7514, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7526, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7556, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7583, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7618, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7652, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7666, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7688, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7709, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7734, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7755, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7764, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7794, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7815, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7808, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7850, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7855, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7859, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7873, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7878, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7900, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7904, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7921, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7929, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7941, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7961, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7967, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7969, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7986, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8003, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8016, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8037, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10697, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13848, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11887, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9467, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8202, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7711, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7562, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7452, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7431, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7444, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7494, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7508, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7553, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7547, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7594, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7612, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7635, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7676, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7684, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7704, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7743, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7740, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7770, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7779, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7803, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7812, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7836, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7840, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7842, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7855, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7876, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7882, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7901, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7927, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7936, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7924, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7965, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7966, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7985, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7995, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8015, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8039, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8074, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10670, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13843, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11905, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9483, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8197, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7722, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7549, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7470, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7439, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7468, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7467, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7503, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7528, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7555, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7580, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7614, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7636, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7656, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7681, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7705, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7735, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7759, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7768, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7779, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7802, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7823, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7825, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7840, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7864, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7880, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7884, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7882, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7905, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7922, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7921, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7952, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7966, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7970, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7980, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7998, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8031, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8038, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8071, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8077, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10637, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13840, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11931, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9495, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8200, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7732, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7544, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7464, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7442, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7446, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7470, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7500, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7526, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7554, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7586, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7628, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7653, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7659, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7687, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7712, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);


	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8073, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8078, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8079, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11054, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13843, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11721, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9367, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8148, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7690, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7545, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7456, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7443, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7439, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7477, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7495, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7518, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7561, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7591, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7636, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7655, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7652, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7700, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7711, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7727, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7749, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7770, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7799, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7780, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7812, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7828, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7841, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7848, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7872, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7887, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7894, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7916, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7919, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7931, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7945, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7959, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7948, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8003, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7998, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8020, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8037, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8076, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11004, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13837, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11735, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9374, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8150, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7696, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7544, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7464, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7439, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7438, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7464, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7502, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7523, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7567, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7596, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7618, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7652, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7662, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7692, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7702, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7742, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7741, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7787, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7788, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7803, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7834, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7835, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7844, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7844, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7867, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7885, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7895, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7901, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7924, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7926, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7944, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7962, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7951, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7982, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8078, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10974, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13831, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11733, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9370, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8157, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7699, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7531, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7472, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7440, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7463, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7471, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7496, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7539, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7547, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7573, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7619, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7648, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7679, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7686, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7722, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7735, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7745, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7787, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7785, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7797, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7818, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7827, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7832, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7864, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7866, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7875, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7899, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7897, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7917, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7934, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7957, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7961, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7980, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7984, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7992, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8016, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8023, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8039, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8034, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8030, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8080, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8079, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10954, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13841, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11766, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9394, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8154, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7696, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7547, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7448, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7427, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7446, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7470, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7504, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7526, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7567, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7596, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7606, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7655, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7665, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7702, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7722, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7730, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7752, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7782, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7777, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7807, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7808, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7839, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7833, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7857, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7862, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7866, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7895, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7909, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7923, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7930, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7942, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7954, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7974, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7979, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7998, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7987, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8016, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8035, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8071, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10900, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13824, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11793, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9403, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8164, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7694, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7544, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7474, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7429, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7436, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7493, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7509, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7540, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7549, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7585, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7613, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7648, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7665, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7695, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7713, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7730, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7746, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7769, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7781, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7812, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7814, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7824, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7840, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7847, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7875, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7876, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7887, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7897, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7909, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7946, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7946, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7965, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7965, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7988, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7997, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8023, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8039, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10866, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13833, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11811, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9422, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8163, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7704, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7548, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7476, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7438, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7452, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7490, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7518, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7534, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7559, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7587, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7631, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7641, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7668, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7685, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7695, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7721, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7760, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7752, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7784, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7816, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7832, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7822, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7843, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7858, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7864, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7876, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7887, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7909, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7907, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7932, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7950, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7949, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7962, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7992, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8007, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8002, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8017, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8037, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10842, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13839, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11810, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9420, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8179, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7711, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7550, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7460, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7438, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7453, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7459, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7486, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7522, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7552, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7570, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7596, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7634, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7672, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7682, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7702, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7727, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7737, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7773, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7796, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7781, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7818, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7830, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7857, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7854, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7865, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7884, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7888, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7898, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7920, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7925, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7945, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7968, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7956, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7999, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8018, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8024, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8032, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8071, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8038, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8041, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10796, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13835, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11838, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9432, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8167, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7708, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7541, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7469, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7442, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7449, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7475, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7508, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7528, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7559, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7575, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7611, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7631, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7654, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7691, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7716, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7722, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7751, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7779, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7791, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7798, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7819, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7829, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7836, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7856, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7872, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7883, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7898, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7903, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7924, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7927, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7950, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7952, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7965, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7973, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8000, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8007, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8034, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8032, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8071, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8076, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8039, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10760, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13837, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11863, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9455, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8172, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7704, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7552, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7476, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7452, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7432, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7484, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7490, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7527, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7564, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7582, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7612, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7636, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7664, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7676, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7710, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7724, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7738, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7763, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7775, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7798, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7821, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7839, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7845, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7857, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7872, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7865, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7884, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7914, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7907, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7926, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7942, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7956, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7967, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7966, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8002, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8004, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8024, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8038, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8035, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8040, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8074, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10749, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13840, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11870, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9461, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8175, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7694, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7548, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7482, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7442, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7434, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7490, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7514, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7526, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7556, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7583, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7618, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7652, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7666, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7688, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7709, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7734, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7755, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7764, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7794, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7815, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7808, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7850, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7855, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7859, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7873, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7878, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7900, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7904, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7921, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7929, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7941, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7961, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7967, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7969, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7986, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8003, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8016, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8037, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8063, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8067, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8045, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8072, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8042, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10697, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13848, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11887, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9467, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8202, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7711, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7562, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7452, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7431, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7444, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7494, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7508, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7553, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7547, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7594, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7612, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7635, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7676, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7684, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7704, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7743, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7740, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7770, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7779, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7803, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7812, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7836, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7840, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7842, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7855, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7876, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7882, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7901, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7927, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7936, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7924, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7965, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7966, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7985, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7995, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8015, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8006, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8039, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8054, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8051, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8052, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8074, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8069, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10670, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13843, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11905, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9483, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8197, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7722, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7549, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7470, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7439, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7468, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7467, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7503, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7528, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7555, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7580, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7614, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7636, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7656, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7681, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7705, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7735, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7759, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7768, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7779, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7802, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7823, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7825, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7840, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7864, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7880, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7884, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7882, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7905, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7922, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7921, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7952, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7966, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7970, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7980, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7998, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8031, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8038, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8066, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8062, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8047, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8064, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8056, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8043, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8060, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8068, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8061, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8055, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8046, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8070, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8057, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8071, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8053, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8059, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8077, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8058, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8049, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8065, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8044, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8048, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8050, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(10637, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(13840, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(11931, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(9495, a2db_data'length);
	a2da_data<=to_unsigned(16383, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(8200, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7732, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7544, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7464, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7442, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7446, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7470, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7500, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7526, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7554, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7586, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7628, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7653, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7659, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7687, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);

	wait for 25 ns;
	a2db_data<=to_unsigned(7712, a2db_data'length);
	a2da_data<=to_unsigned(0, a2da_data'length);


				
		
		
	end process;
	
		
		
end behave;