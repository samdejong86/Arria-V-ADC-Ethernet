-- Nios_CPU_qsys.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Nios_CPU_qsys is
	port (
		adc_control_out_export                          : out   std_logic_vector(7 downto 0);                     --                     adc_control_out.export
		cfi_flash_atb_bridge_0_out_tcm_address_out      : out   std_logic_vector(26 downto 0);                    --          cfi_flash_atb_bridge_0_out.tcm_address_out
		cfi_flash_atb_bridge_0_out_tcm_read_n_out       : out   std_logic_vector(0 downto 0);                     --                                    .tcm_read_n_out
		cfi_flash_atb_bridge_0_out_tcm_write_n_out      : out   std_logic_vector(0 downto 0);                     --                                    .tcm_write_n_out
		cfi_flash_atb_bridge_0_out_tcm_data_out         : inout std_logic_vector(15 downto 0) := (others => '0'); --                                    .tcm_data_out
		cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out : out   std_logic_vector(0 downto 0);                     --                                    .tcm_chipselect_n_out
		clk_clk                                         : in    std_logic                     := '0';             --                                 clk.clk
		enet_pll_locked_export                          : out   std_logic;                                        --                     enet_pll_locked.export
		enet_pll_outclk0_clk                            : out   std_logic;                                        --                    enet_pll_outclk0.clk
		enet_pll_outclk1_clk                            : out   std_logic;                                        --                    enet_pll_outclk1.clk
		enet_pll_outclk2_clk                            : out   std_logic;                                        --                    enet_pll_outclk2.clk
		enet_pll_reset_reset                            : in    std_logic                     := '0';             --                      enet_pll_reset.reset
		lcd_external_RS                                 : out   std_logic;                                        --                        lcd_external.RS
		lcd_external_RW                                 : out   std_logic;                                        --                                    .RW
		lcd_external_data                               : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                    .data
		lcd_external_E                                  : out   std_logic;                                        --                                    .E
		merged_resets_in_reset_reset_n                  : in    std_logic                     := '0';             --              merged_resets_in_reset.reset_n
		samplenum_out_export                            : out   std_logic_vector(15 downto 0);                    --                       samplenum_out.export
		tse_mac_mac_mdio_connection_mdc                 : out   std_logic;                                        --         tse_mac_mac_mdio_connection.mdc
		tse_mac_mac_mdio_connection_mdio_in             : in    std_logic                     := '0';             --                                    .mdio_in
		tse_mac_mac_mdio_connection_mdio_out            : out   std_logic;                                        --                                    .mdio_out
		tse_mac_mac_mdio_connection_mdio_oen            : out   std_logic;                                        --                                    .mdio_oen
		tse_mac_mac_rgmii_connection_rgmii_in           : in    std_logic_vector(3 downto 0)  := (others => '0'); --        tse_mac_mac_rgmii_connection.rgmii_in
		tse_mac_mac_rgmii_connection_rgmii_out          : out   std_logic_vector(3 downto 0);                     --                                    .rgmii_out
		tse_mac_mac_rgmii_connection_rx_control         : in    std_logic                     := '0';             --                                    .rx_control
		tse_mac_mac_rgmii_connection_tx_control         : out   std_logic;                                        --                                    .tx_control
		tse_mac_mac_status_connection_set_10            : in    std_logic                     := '0';             --       tse_mac_mac_status_connection.set_10
		tse_mac_mac_status_connection_set_1000          : in    std_logic                     := '0';             --                                    .set_1000
		tse_mac_mac_status_connection_eth_mode          : out   std_logic;                                        --                                    .eth_mode
		tse_mac_mac_status_connection_ena_10            : out   std_logic;                                        --                                    .ena_10
		tse_mac_pcs_mac_rx_clock_connection_clk         : in    std_logic                     := '0';             -- tse_mac_pcs_mac_rx_clock_connection.clk
		tse_mac_pcs_mac_tx_clock_connection_clk         : in    std_logic                     := '0';             -- tse_mac_pcs_mac_tx_clock_connection.clk
		wavesample_in_export                            : in    std_logic_vector(15 downto 0) := (others => '0')  --                       wavesample_in.export
	);
end entity Nios_CPU_qsys;

architecture rtl of Nios_CPU_qsys is
	component Nios_CPU_qsys_adc_control is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component Nios_CPU_qsys_adc_control;

	component Nios_CPU_qsys_cfi_flash_atb_bridge_0 is
		port (
			clk                      : in    std_logic                     := 'X';             -- clk
			reset                    : in    std_logic                     := 'X';             -- reset
			request                  : in    std_logic                     := 'X';             -- request
			grant                    : out   std_logic;                                        -- grant
			tcs_tcm_address_out      : in    std_logic_vector(26 downto 0) := (others => 'X'); -- address_out
			tcs_tcm_read_n_out       : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- read_n_out
			tcs_tcm_write_n_out      : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_out
			tcs_tcm_data_out         : in    std_logic_vector(15 downto 0) := (others => 'X'); -- data_out
			tcs_tcm_data_outen       : in    std_logic                     := 'X';             -- data_outen
			tcs_tcm_data_in          : out   std_logic_vector(15 downto 0);                    -- data_in
			tcs_tcm_chipselect_n_out : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- chipselect_n_out
			tcm_address_out          : out   std_logic_vector(26 downto 0);                    -- tcm_address_out
			tcm_read_n_out           : out   std_logic_vector(0 downto 0);                     -- tcm_read_n_out
			tcm_write_n_out          : out   std_logic_vector(0 downto 0);                     -- tcm_write_n_out
			tcm_data_out             : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			tcm_chipselect_n_out     : out   std_logic_vector(0 downto 0)                      -- tcm_chipselect_n_out
		);
	end component Nios_CPU_qsys_cfi_flash_atb_bridge_0;

	component Nios_CPU_qsys_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component Nios_CPU_qsys_cpu;

	component Nios_CPU_qsys_descriptor_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component Nios_CPU_qsys_descriptor_memory;

	component Nios_CPU_qsys_enet_pll is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component Nios_CPU_qsys_enet_pll;

	component Nios_CPU_qsys_ext_flash is
		generic (
			TCM_ADDRESS_W                  : integer := 30;
			TCM_DATA_W                     : integer := 32;
			TCM_BYTEENABLE_W               : integer := 4;
			TCM_READ_WAIT                  : integer := 1;
			TCM_WRITE_WAIT                 : integer := 0;
			TCM_SETUP_WAIT                 : integer := 0;
			TCM_DATA_HOLD                  : integer := 0;
			TCM_TURNAROUND_TIME            : integer := 2;
			TCM_TIMING_UNITS               : integer := 1;
			TCM_READLATENCY                : integer := 2;
			TCM_SYMBOLS_PER_WORD           : integer := 4;
			USE_READDATA                   : integer := 1;
			USE_WRITEDATA                  : integer := 1;
			USE_READ                       : integer := 1;
			USE_WRITE                      : integer := 1;
			USE_BYTEENABLE                 : integer := 1;
			USE_CHIPSELECT                 : integer := 0;
			USE_LOCK                       : integer := 0;
			USE_ADDRESS                    : integer := 1;
			USE_WAITREQUEST                : integer := 0;
			USE_WRITEBYTEENABLE            : integer := 0;
			USE_OUTPUTENABLE               : integer := 0;
			USE_RESETREQUEST               : integer := 0;
			USE_IRQ                        : integer := 0;
			USE_RESET_OUTPUT               : integer := 0;
			ACTIVE_LOW_READ                : integer := 0;
			ACTIVE_LOW_LOCK                : integer := 0;
			ACTIVE_LOW_WRITE               : integer := 0;
			ACTIVE_LOW_CHIPSELECT          : integer := 0;
			ACTIVE_LOW_BYTEENABLE          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE        : integer := 0;
			ACTIVE_LOW_WRITEBYTEENABLE     : integer := 0;
			ACTIVE_LOW_WAITREQUEST         : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER       : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			reset_reset          : in  std_logic                     := 'X';             -- reset
			uas_address          : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			uas_burstcount       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uas_read             : in  std_logic                     := 'X';             -- read
			uas_write            : in  std_logic                     := 'X';             -- write
			uas_waitrequest      : out std_logic;                                        -- waitrequest
			uas_readdatavalid    : out std_logic;                                        -- readdatavalid
			uas_byteenable       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uas_readdata         : out std_logic_vector(15 downto 0);                    -- readdata
			uas_writedata        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uas_lock             : in  std_logic                     := 'X';             -- lock
			uas_debugaccess      : in  std_logic                     := 'X';             -- debugaccess
			tcm_write_n_out      : out std_logic;                                        -- write_n_out
			tcm_read_n_out       : out std_logic;                                        -- read_n_out
			tcm_chipselect_n_out : out std_logic;                                        -- chipselect_n_out
			tcm_request          : out std_logic;                                        -- request
			tcm_grant            : in  std_logic                     := 'X';             -- grant
			tcm_address_out      : out std_logic_vector(26 downto 0);                    -- address_out
			tcm_data_out         : out std_logic_vector(15 downto 0);                    -- data_out
			tcm_data_outen       : out std_logic;                                        -- data_outen
			tcm_data_in          : in  std_logic_vector(15 downto 0) := (others => 'X')  -- data_in
		);
	end component Nios_CPU_qsys_ext_flash;

	component Nios_CPU_qsys_high_res_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component Nios_CPU_qsys_high_res_timer;

	component Nios_CPU_qsys_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Nios_CPU_qsys_jtag_uart_0;

	component Nios_CPU_qsys_lcd is
		port (
			reset_n       : in    std_logic                    := 'X';             -- reset_n
			clk           : in    std_logic                    := 'X';             -- clk
			begintransfer : in    std_logic                    := 'X';             -- begintransfer
			read          : in    std_logic                    := 'X';             -- read
			write         : in    std_logic                    := 'X';             -- write
			readdata      : out   std_logic_vector(7 downto 0);                    -- readdata
			writedata     : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			address       : in    std_logic_vector(1 downto 0) := (others => 'X'); -- address
			LCD_RS        : out   std_logic;                                       -- export
			LCD_RW        : out   std_logic;                                       -- export
			LCD_data      : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			LCD_E         : out   std_logic                                        -- export
		);
	end component Nios_CPU_qsys_lcd;

	component Nios_CPU_qsys_onchip_ram is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component Nios_CPU_qsys_onchip_ram;

	component altera_avalon_mm_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(9 downto 0);                     -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component altera_avalon_mm_bridge;

	component Nios_CPU_qsys_sampleNum is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(15 downto 0)                     -- export
		);
	end component Nios_CPU_qsys_sampleNum;

	component Nios_CPU_qsys_sgdma_rx is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			in_startofpacket              : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket                : in  std_logic                     := 'X';             -- endofpacket
			in_data                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_valid                      : in  std_logic                     := 'X';             -- valid
			in_ready                      : out std_logic;                                        -- ready
			in_empty                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			in_error                      : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- error
			m_write_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			m_write_address               : out std_logic_vector(31 downto 0);                    -- address
			m_write_write                 : out std_logic;                                        -- write
			m_write_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			m_write_byteenable            : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component Nios_CPU_qsys_sgdma_rx;

	component Nios_CPU_qsys_sgdma_tx is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			m_read_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m_read_readdatavalid          : in  std_logic                     := 'X';             -- readdatavalid
			m_read_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			m_read_address                : out std_logic_vector(31 downto 0);                    -- address
			m_read_read                   : out std_logic;                                        -- read
			out_data                      : out std_logic_vector(31 downto 0);                    -- data
			out_valid                     : out std_logic;                                        -- valid
			out_ready                     : in  std_logic                     := 'X';             -- ready
			out_endofpacket               : out std_logic;                                        -- endofpacket
			out_startofpacket             : out std_logic;                                        -- startofpacket
			out_empty                     : out std_logic_vector(1 downto 0);                     -- empty
			out_error                     : out std_logic                                         -- error
		);
	end component Nios_CPU_qsys_sgdma_tx;

	component Nios_CPU_qsys_sys_clk_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component Nios_CPU_qsys_sys_clk_timer;

	component Nios_CPU_qsys_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component Nios_CPU_qsys_sysid;

	component Nios_CPU_qsys_tse_mac is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			reg_addr      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			reg_data_out  : out std_logic_vector(31 downto 0);                    -- readdata
			reg_rd        : in  std_logic                     := 'X';             -- read
			reg_data_in   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reg_wr        : in  std_logic                     := 'X';             -- write
			reg_busy      : out std_logic;                                        -- waitrequest
			tx_clk        : in  std_logic                     := 'X';             -- clk
			rx_clk        : in  std_logic                     := 'X';             -- clk
			set_10        : in  std_logic                     := 'X';             -- set_10
			set_1000      : in  std_logic                     := 'X';             -- set_1000
			eth_mode      : out std_logic;                                        -- eth_mode
			ena_10        : out std_logic;                                        -- ena_10
			rgmii_in      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- rgmii_in
			rgmii_out     : out std_logic_vector(3 downto 0);                     -- rgmii_out
			rx_control    : in  std_logic                     := 'X';             -- rx_control
			tx_control    : out std_logic;                                        -- tx_control
			ff_rx_clk     : in  std_logic                     := 'X';             -- clk
			ff_tx_clk     : in  std_logic                     := 'X';             -- clk
			ff_rx_data    : out std_logic_vector(31 downto 0);                    -- data
			ff_rx_eop     : out std_logic;                                        -- endofpacket
			rx_err        : out std_logic_vector(5 downto 0);                     -- error
			ff_rx_mod     : out std_logic_vector(1 downto 0);                     -- empty
			ff_rx_rdy     : in  std_logic                     := 'X';             -- ready
			ff_rx_sop     : out std_logic;                                        -- startofpacket
			ff_rx_dval    : out std_logic;                                        -- valid
			ff_tx_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			ff_tx_eop     : in  std_logic                     := 'X';             -- endofpacket
			ff_tx_err     : in  std_logic                     := 'X';             -- error
			ff_tx_mod     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			ff_tx_rdy     : out std_logic;                                        -- ready
			ff_tx_sop     : in  std_logic                     := 'X';             -- startofpacket
			ff_tx_wren    : in  std_logic                     := 'X';             -- valid
			mdc           : out std_logic;                                        -- mdc
			mdio_in       : in  std_logic                     := 'X';             -- mdio_in
			mdio_out      : out std_logic;                                        -- mdio_out
			mdio_oen      : out std_logic;                                        -- mdio_oen
			xon_gen       : in  std_logic                     := 'X';             -- xon_gen
			xoff_gen      : in  std_logic                     := 'X';             -- xoff_gen
			ff_tx_crc_fwd : in  std_logic                     := 'X';             -- ff_tx_crc_fwd
			ff_tx_septy   : out std_logic;                                        -- ff_tx_septy
			tx_ff_uflow   : out std_logic;                                        -- tx_ff_uflow
			ff_tx_a_full  : out std_logic;                                        -- ff_tx_a_full
			ff_tx_a_empty : out std_logic;                                        -- ff_tx_a_empty
			rx_err_stat   : out std_logic_vector(17 downto 0);                    -- rx_err_stat
			rx_frm_type   : out std_logic_vector(3 downto 0);                     -- rx_frm_type
			ff_rx_dsav    : out std_logic;                                        -- ff_rx_dsav
			ff_rx_a_full  : out std_logic;                                        -- ff_rx_a_full
			ff_rx_a_empty : out std_logic                                         -- ff_rx_a_empty
		);
	end component Nios_CPU_qsys_tse_mac;

	component Nios_CPU_qsys_waveSample is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(15 downto 0) := (others => 'X')  -- export
		);
	end component Nios_CPU_qsys_waveSample;

	component Nios_CPU_qsys_mm_interconnect_0 is
		port (
			clkin_50_clk_clk                           : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset      : in  std_logic                     := 'X';             -- reset
			sgdma_tx_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                    : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                       : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_readdatavalid              : out std_logic;                                        -- readdatavalid
			cpu_data_master_write                      : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address             : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest         : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_instruction_master_readdatavalid       : out std_logic;                                        -- readdatavalid
			sgdma_rx_descriptor_read_address           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_rx_descriptor_read_waitrequest       : out std_logic;                                        -- waitrequest
			sgdma_rx_descriptor_read_read              : in  std_logic                     := 'X';             -- read
			sgdma_rx_descriptor_read_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			sgdma_rx_descriptor_read_readdatavalid     : out std_logic;                                        -- readdatavalid
			sgdma_rx_descriptor_write_address          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_rx_descriptor_write_waitrequest      : out std_logic;                                        -- waitrequest
			sgdma_rx_descriptor_write_write            : in  std_logic                     := 'X';             -- write
			sgdma_rx_descriptor_write_writedata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sgdma_rx_m_write_address                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_rx_m_write_waitrequest               : out std_logic;                                        -- waitrequest
			sgdma_rx_m_write_byteenable                : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			sgdma_rx_m_write_write                     : in  std_logic                     := 'X';             -- write
			sgdma_rx_m_write_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sgdma_tx_descriptor_read_address           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_tx_descriptor_read_waitrequest       : out std_logic;                                        -- waitrequest
			sgdma_tx_descriptor_read_read              : in  std_logic                     := 'X';             -- read
			sgdma_tx_descriptor_read_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			sgdma_tx_descriptor_read_readdatavalid     : out std_logic;                                        -- readdatavalid
			sgdma_tx_descriptor_write_address          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_tx_descriptor_write_waitrequest      : out std_logic;                                        -- waitrequest
			sgdma_tx_descriptor_write_write            : in  std_logic                     := 'X';             -- write
			sgdma_tx_descriptor_write_writedata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sgdma_tx_m_read_address                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_tx_m_read_waitrequest                : out std_logic;                                        -- waitrequest
			sgdma_tx_m_read_read                       : in  std_logic                     := 'X';             -- read
			sgdma_tx_m_read_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			sgdma_tx_m_read_readdatavalid              : out std_logic;                                        -- readdatavalid
			cpu_debug_mem_slave_address                : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                  : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                   : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable             : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess            : out std_logic;                                        -- debugaccess
			descriptor_memory_s1_address               : out std_logic_vector(10 downto 0);                    -- address
			descriptor_memory_s1_write                 : out std_logic;                                        -- write
			descriptor_memory_s1_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_memory_s1_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			descriptor_memory_s1_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			descriptor_memory_s1_chipselect            : out std_logic;                                        -- chipselect
			descriptor_memory_s1_clken                 : out std_logic;                                        -- clken
			ext_flash_uas_address                      : out std_logic_vector(26 downto 0);                    -- address
			ext_flash_uas_write                        : out std_logic;                                        -- write
			ext_flash_uas_read                         : out std_logic;                                        -- read
			ext_flash_uas_readdata                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			ext_flash_uas_writedata                    : out std_logic_vector(15 downto 0);                    -- writedata
			ext_flash_uas_burstcount                   : out std_logic_vector(1 downto 0);                     -- burstcount
			ext_flash_uas_byteenable                   : out std_logic_vector(1 downto 0);                     -- byteenable
			ext_flash_uas_readdatavalid                : in  std_logic                     := 'X';             -- readdatavalid
			ext_flash_uas_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			ext_flash_uas_lock                         : out std_logic;                                        -- lock
			ext_flash_uas_debugaccess                  : out std_logic;                                        -- debugaccess
			onchip_ram_s1_address                      : out std_logic_vector(18 downto 0);                    -- address
			onchip_ram_s1_write                        : out std_logic;                                        -- write
			onchip_ram_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_ram_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_ram_s1_byteenable                   : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_ram_s1_chipselect                   : out std_logic;                                        -- chipselect
			onchip_ram_s1_clken                        : out std_logic;                                        -- clken
			onchip_ram_s2_address                      : out std_logic_vector(18 downto 0);                    -- address
			onchip_ram_s2_write                        : out std_logic;                                        -- write
			onchip_ram_s2_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_ram_s2_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_ram_s2_byteenable                   : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_ram_s2_chipselect                   : out std_logic;                                        -- chipselect
			onchip_ram_s2_clken                        : out std_logic;                                        -- clken
			pb_cpu_to_io_s0_address                    : out std_logic_vector(9 downto 0);                     -- address
			pb_cpu_to_io_s0_write                      : out std_logic;                                        -- write
			pb_cpu_to_io_s0_read                       : out std_logic;                                        -- read
			pb_cpu_to_io_s0_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pb_cpu_to_io_s0_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			pb_cpu_to_io_s0_burstcount                 : out std_logic_vector(0 downto 0);                     -- burstcount
			pb_cpu_to_io_s0_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			pb_cpu_to_io_s0_readdatavalid              : in  std_logic                     := 'X';             -- readdatavalid
			pb_cpu_to_io_s0_waitrequest                : in  std_logic                     := 'X';             -- waitrequest
			pb_cpu_to_io_s0_debugaccess                : out std_logic;                                        -- debugaccess
			sgdma_rx_csr_address                       : out std_logic_vector(3 downto 0);                     -- address
			sgdma_rx_csr_write                         : out std_logic;                                        -- write
			sgdma_rx_csr_read                          : out std_logic;                                        -- read
			sgdma_rx_csr_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sgdma_rx_csr_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			sgdma_rx_csr_chipselect                    : out std_logic;                                        -- chipselect
			sgdma_tx_csr_address                       : out std_logic_vector(3 downto 0);                     -- address
			sgdma_tx_csr_write                         : out std_logic;                                        -- write
			sgdma_tx_csr_read                          : out std_logic;                                        -- read
			sgdma_tx_csr_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sgdma_tx_csr_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			sgdma_tx_csr_chipselect                    : out std_logic;                                        -- chipselect
			tse_mac_control_port_address               : out std_logic_vector(7 downto 0);                     -- address
			tse_mac_control_port_write                 : out std_logic;                                        -- write
			tse_mac_control_port_read                  : out std_logic;                                        -- read
			tse_mac_control_port_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			tse_mac_control_port_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			tse_mac_control_port_waitrequest           : in  std_logic                     := 'X'              -- waitrequest
		);
	end component Nios_CPU_qsys_mm_interconnect_0;

	component Nios_CPU_qsys_mm_interconnect_1 is
		port (
			clkin_50_clk_clk                               : in  std_logic                     := 'X';             -- clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			pb_cpu_to_io_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			pb_cpu_to_io_m0_address                        : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			pb_cpu_to_io_m0_waitrequest                    : out std_logic;                                        -- waitrequest
			pb_cpu_to_io_m0_burstcount                     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			pb_cpu_to_io_m0_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			pb_cpu_to_io_m0_read                           : in  std_logic                     := 'X';             -- read
			pb_cpu_to_io_m0_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			pb_cpu_to_io_m0_readdatavalid                  : out std_logic;                                        -- readdatavalid
			pb_cpu_to_io_m0_write                          : in  std_logic                     := 'X';             -- write
			pb_cpu_to_io_m0_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pb_cpu_to_io_m0_debugaccess                    : in  std_logic                     := 'X';             -- debugaccess
			adc_control_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			adc_control_s1_write                           : out std_logic;                                        -- write
			adc_control_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			adc_control_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			adc_control_s1_chipselect                      : out std_logic;                                        -- chipselect
			high_res_timer_s1_address                      : out std_logic_vector(2 downto 0);                     -- address
			high_res_timer_s1_write                        : out std_logic;                                        -- write
			high_res_timer_s1_readdata                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			high_res_timer_s1_writedata                    : out std_logic_vector(15 downto 0);                    -- writedata
			high_res_timer_s1_chipselect                   : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address          : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write            : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read             : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect       : out std_logic;                                        -- chipselect
			lcd_control_slave_address                      : out std_logic_vector(1 downto 0);                     -- address
			lcd_control_slave_write                        : out std_logic;                                        -- write
			lcd_control_slave_read                         : out std_logic;                                        -- read
			lcd_control_slave_readdata                     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			lcd_control_slave_writedata                    : out std_logic_vector(7 downto 0);                     -- writedata
			lcd_control_slave_begintransfer                : out std_logic;                                        -- begintransfer
			sampleNum_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			sampleNum_s1_write                             : out std_logic;                                        -- write
			sampleNum_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sampleNum_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			sampleNum_s1_chipselect                        : out std_logic;                                        -- chipselect
			sys_clk_timer_s1_address                       : out std_logic_vector(2 downto 0);                     -- address
			sys_clk_timer_s1_write                         : out std_logic;                                        -- write
			sys_clk_timer_s1_readdata                      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sys_clk_timer_s1_writedata                     : out std_logic_vector(15 downto 0);                    -- writedata
			sys_clk_timer_s1_chipselect                    : out std_logic;                                        -- chipselect
			sysid_control_slave_address                    : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			waveSample_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			waveSample_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component Nios_CPU_qsys_mm_interconnect_1;

	component Nios_CPU_qsys_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Nios_CPU_qsys_irq_mapper;

	component Nios_CPU_qsys_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_empty          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			in_0_error          : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- error
			out_0_data          : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic;                                        -- endofpacket
			out_0_empty         : out std_logic_vector(1 downto 0);                     -- empty
			out_0_error         : out std_logic_vector(5 downto 0)                      -- error
		);
	end component Nios_CPU_qsys_avalon_st_adapter;

	component nios_cpu_qsys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_cpu_qsys_rst_controller;

	component nios_cpu_qsys_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_in2      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_cpu_qsys_rst_controller_001;

	signal sgdma_tx_out_valid                                              : std_logic;                     -- sgdma_tx:out_valid -> tse_mac:ff_tx_wren
	signal sgdma_tx_out_data                                               : std_logic_vector(31 downto 0); -- sgdma_tx:out_data -> tse_mac:ff_tx_data
	signal sgdma_tx_out_ready                                              : std_logic;                     -- tse_mac:ff_tx_rdy -> sgdma_tx:out_ready
	signal sgdma_tx_out_startofpacket                                      : std_logic;                     -- sgdma_tx:out_startofpacket -> tse_mac:ff_tx_sop
	signal sgdma_tx_out_endofpacket                                        : std_logic;                     -- sgdma_tx:out_endofpacket -> tse_mac:ff_tx_eop
	signal sgdma_tx_out_error                                              : std_logic;                     -- sgdma_tx:out_error -> tse_mac:ff_tx_err
	signal sgdma_tx_out_empty                                              : std_logic_vector(1 downto 0);  -- sgdma_tx:out_empty -> tse_mac:ff_tx_mod
	signal ext_flash_tcm_data_outen                                        : std_logic;                     -- ext_flash:tcm_data_outen -> cfi_flash_atb_bridge_0:tcs_tcm_data_outen
	signal ext_flash_tcm_request                                           : std_logic;                     -- ext_flash:tcm_request -> cfi_flash_atb_bridge_0:request
	signal ext_flash_tcm_write_n_out                                       : std_logic;                     -- ext_flash:tcm_write_n_out -> cfi_flash_atb_bridge_0:tcs_tcm_write_n_out
	signal ext_flash_tcm_read_n_out                                        : std_logic;                     -- ext_flash:tcm_read_n_out -> cfi_flash_atb_bridge_0:tcs_tcm_read_n_out
	signal ext_flash_tcm_grant                                             : std_logic;                     -- cfi_flash_atb_bridge_0:grant -> ext_flash:tcm_grant
	signal ext_flash_tcm_chipselect_n_out                                  : std_logic;                     -- ext_flash:tcm_chipselect_n_out -> cfi_flash_atb_bridge_0:tcs_tcm_chipselect_n_out
	signal ext_flash_tcm_address_out                                       : std_logic_vector(26 downto 0); -- ext_flash:tcm_address_out -> cfi_flash_atb_bridge_0:tcs_tcm_address_out
	signal ext_flash_tcm_data_out                                          : std_logic_vector(15 downto 0); -- ext_flash:tcm_data_out -> cfi_flash_atb_bridge_0:tcs_tcm_data_out
	signal ext_flash_tcm_data_in                                           : std_logic_vector(15 downto 0); -- cfi_flash_atb_bridge_0:tcs_tcm_data_in -> ext_flash:tcm_data_in
	signal cpu_data_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                     : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                         : std_logic_vector(27 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                      : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                            : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	signal cpu_data_master_write                                           : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                       : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                  : std_logic_vector(27 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                     : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal cpu_instruction_master_readdatavalid                            : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	signal sgdma_tx_m_read_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_tx_m_read_readdata -> sgdma_tx:m_read_readdata
	signal sgdma_tx_m_read_waitrequest                                     : std_logic;                     -- mm_interconnect_0:sgdma_tx_m_read_waitrequest -> sgdma_tx:m_read_waitrequest
	signal sgdma_tx_m_read_address                                         : std_logic_vector(31 downto 0); -- sgdma_tx:m_read_address -> mm_interconnect_0:sgdma_tx_m_read_address
	signal sgdma_tx_m_read_read                                            : std_logic;                     -- sgdma_tx:m_read_read -> mm_interconnect_0:sgdma_tx_m_read_read
	signal sgdma_tx_m_read_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:sgdma_tx_m_read_readdatavalid -> sgdma_tx:m_read_readdatavalid
	signal sgdma_rx_m_write_waitrequest                                    : std_logic;                     -- mm_interconnect_0:sgdma_rx_m_write_waitrequest -> sgdma_rx:m_write_waitrequest
	signal sgdma_rx_m_write_address                                        : std_logic_vector(31 downto 0); -- sgdma_rx:m_write_address -> mm_interconnect_0:sgdma_rx_m_write_address
	signal sgdma_rx_m_write_byteenable                                     : std_logic_vector(3 downto 0);  -- sgdma_rx:m_write_byteenable -> mm_interconnect_0:sgdma_rx_m_write_byteenable
	signal sgdma_rx_m_write_write                                          : std_logic;                     -- sgdma_rx:m_write_write -> mm_interconnect_0:sgdma_rx_m_write_write
	signal sgdma_rx_m_write_writedata                                      : std_logic_vector(31 downto 0); -- sgdma_rx:m_write_writedata -> mm_interconnect_0:sgdma_rx_m_write_writedata
	signal sgdma_rx_descriptor_read_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_rx_descriptor_read_readdata -> sgdma_rx:descriptor_read_readdata
	signal sgdma_rx_descriptor_read_waitrequest                            : std_logic;                     -- mm_interconnect_0:sgdma_rx_descriptor_read_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	signal sgdma_rx_descriptor_read_address                                : std_logic_vector(31 downto 0); -- sgdma_rx:descriptor_read_address -> mm_interconnect_0:sgdma_rx_descriptor_read_address
	signal sgdma_rx_descriptor_read_read                                   : std_logic;                     -- sgdma_rx:descriptor_read_read -> mm_interconnect_0:sgdma_rx_descriptor_read_read
	signal sgdma_rx_descriptor_read_readdatavalid                          : std_logic;                     -- mm_interconnect_0:sgdma_rx_descriptor_read_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	signal sgdma_tx_descriptor_read_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_tx_descriptor_read_readdata -> sgdma_tx:descriptor_read_readdata
	signal sgdma_tx_descriptor_read_waitrequest                            : std_logic;                     -- mm_interconnect_0:sgdma_tx_descriptor_read_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	signal sgdma_tx_descriptor_read_address                                : std_logic_vector(31 downto 0); -- sgdma_tx:descriptor_read_address -> mm_interconnect_0:sgdma_tx_descriptor_read_address
	signal sgdma_tx_descriptor_read_read                                   : std_logic;                     -- sgdma_tx:descriptor_read_read -> mm_interconnect_0:sgdma_tx_descriptor_read_read
	signal sgdma_tx_descriptor_read_readdatavalid                          : std_logic;                     -- mm_interconnect_0:sgdma_tx_descriptor_read_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	signal sgdma_rx_descriptor_write_waitrequest                           : std_logic;                     -- mm_interconnect_0:sgdma_rx_descriptor_write_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	signal sgdma_rx_descriptor_write_address                               : std_logic_vector(31 downto 0); -- sgdma_rx:descriptor_write_address -> mm_interconnect_0:sgdma_rx_descriptor_write_address
	signal sgdma_rx_descriptor_write_write                                 : std_logic;                     -- sgdma_rx:descriptor_write_write -> mm_interconnect_0:sgdma_rx_descriptor_write_write
	signal sgdma_rx_descriptor_write_writedata                             : std_logic_vector(31 downto 0); -- sgdma_rx:descriptor_write_writedata -> mm_interconnect_0:sgdma_rx_descriptor_write_writedata
	signal sgdma_tx_descriptor_write_waitrequest                           : std_logic;                     -- mm_interconnect_0:sgdma_tx_descriptor_write_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	signal sgdma_tx_descriptor_write_address                               : std_logic_vector(31 downto 0); -- sgdma_tx:descriptor_write_address -> mm_interconnect_0:sgdma_tx_descriptor_write_address
	signal sgdma_tx_descriptor_write_write                                 : std_logic;                     -- sgdma_tx:descriptor_write_write -> mm_interconnect_0:sgdma_tx_descriptor_write_write
	signal sgdma_tx_descriptor_write_writedata                             : std_logic_vector(31 downto 0); -- sgdma_tx:descriptor_write_writedata -> mm_interconnect_0:sgdma_tx_descriptor_write_writedata
	signal mm_interconnect_0_tse_mac_control_port_readdata                 : std_logic_vector(31 downto 0); -- tse_mac:reg_data_out -> mm_interconnect_0:tse_mac_control_port_readdata
	signal mm_interconnect_0_tse_mac_control_port_waitrequest              : std_logic;                     -- tse_mac:reg_busy -> mm_interconnect_0:tse_mac_control_port_waitrequest
	signal mm_interconnect_0_tse_mac_control_port_address                  : std_logic_vector(7 downto 0);  -- mm_interconnect_0:tse_mac_control_port_address -> tse_mac:reg_addr
	signal mm_interconnect_0_tse_mac_control_port_read                     : std_logic;                     -- mm_interconnect_0:tse_mac_control_port_read -> tse_mac:reg_rd
	signal mm_interconnect_0_tse_mac_control_port_write                    : std_logic;                     -- mm_interconnect_0:tse_mac_control_port_write -> tse_mac:reg_wr
	signal mm_interconnect_0_tse_mac_control_port_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:tse_mac_control_port_writedata -> tse_mac:reg_data_in
	signal mm_interconnect_0_sgdma_tx_csr_chipselect                       : std_logic;                     -- mm_interconnect_0:sgdma_tx_csr_chipselect -> sgdma_tx:csr_chipselect
	signal mm_interconnect_0_sgdma_tx_csr_readdata                         : std_logic_vector(31 downto 0); -- sgdma_tx:csr_readdata -> mm_interconnect_0:sgdma_tx_csr_readdata
	signal mm_interconnect_0_sgdma_tx_csr_address                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sgdma_tx_csr_address -> sgdma_tx:csr_address
	signal mm_interconnect_0_sgdma_tx_csr_read                             : std_logic;                     -- mm_interconnect_0:sgdma_tx_csr_read -> sgdma_tx:csr_read
	signal mm_interconnect_0_sgdma_tx_csr_write                            : std_logic;                     -- mm_interconnect_0:sgdma_tx_csr_write -> sgdma_tx:csr_write
	signal mm_interconnect_0_sgdma_tx_csr_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_tx_csr_writedata -> sgdma_tx:csr_writedata
	signal mm_interconnect_0_sgdma_rx_csr_chipselect                       : std_logic;                     -- mm_interconnect_0:sgdma_rx_csr_chipselect -> sgdma_rx:csr_chipselect
	signal mm_interconnect_0_sgdma_rx_csr_readdata                         : std_logic_vector(31 downto 0); -- sgdma_rx:csr_readdata -> mm_interconnect_0:sgdma_rx_csr_readdata
	signal mm_interconnect_0_sgdma_rx_csr_address                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sgdma_rx_csr_address -> sgdma_rx:csr_address
	signal mm_interconnect_0_sgdma_rx_csr_read                             : std_logic;                     -- mm_interconnect_0:sgdma_rx_csr_read -> sgdma_rx:csr_read
	signal mm_interconnect_0_sgdma_rx_csr_write                            : std_logic;                     -- mm_interconnect_0:sgdma_rx_csr_write -> sgdma_rx:csr_write
	signal mm_interconnect_0_sgdma_rx_csr_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_rx_csr_writedata -> sgdma_rx:csr_writedata
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                  : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest               : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess               : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                   : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                      : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                     : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_pb_cpu_to_io_s0_readdata                      : std_logic_vector(31 downto 0); -- pb_cpu_to_io:s0_readdata -> mm_interconnect_0:pb_cpu_to_io_s0_readdata
	signal mm_interconnect_0_pb_cpu_to_io_s0_waitrequest                   : std_logic;                     -- pb_cpu_to_io:s0_waitrequest -> mm_interconnect_0:pb_cpu_to_io_s0_waitrequest
	signal mm_interconnect_0_pb_cpu_to_io_s0_debugaccess                   : std_logic;                     -- mm_interconnect_0:pb_cpu_to_io_s0_debugaccess -> pb_cpu_to_io:s0_debugaccess
	signal mm_interconnect_0_pb_cpu_to_io_s0_address                       : std_logic_vector(9 downto 0);  -- mm_interconnect_0:pb_cpu_to_io_s0_address -> pb_cpu_to_io:s0_address
	signal mm_interconnect_0_pb_cpu_to_io_s0_read                          : std_logic;                     -- mm_interconnect_0:pb_cpu_to_io_s0_read -> pb_cpu_to_io:s0_read
	signal mm_interconnect_0_pb_cpu_to_io_s0_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:pb_cpu_to_io_s0_byteenable -> pb_cpu_to_io:s0_byteenable
	signal mm_interconnect_0_pb_cpu_to_io_s0_readdatavalid                 : std_logic;                     -- pb_cpu_to_io:s0_readdatavalid -> mm_interconnect_0:pb_cpu_to_io_s0_readdatavalid
	signal mm_interconnect_0_pb_cpu_to_io_s0_write                         : std_logic;                     -- mm_interconnect_0:pb_cpu_to_io_s0_write -> pb_cpu_to_io:s0_write
	signal mm_interconnect_0_pb_cpu_to_io_s0_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:pb_cpu_to_io_s0_writedata -> pb_cpu_to_io:s0_writedata
	signal mm_interconnect_0_pb_cpu_to_io_s0_burstcount                    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:pb_cpu_to_io_s0_burstcount -> pb_cpu_to_io:s0_burstcount
	signal mm_interconnect_0_onchip_ram_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	signal mm_interconnect_0_onchip_ram_s1_readdata                        : std_logic_vector(31 downto 0); -- onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	signal mm_interconnect_0_onchip_ram_s1_address                         : std_logic_vector(18 downto 0); -- mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	signal mm_interconnect_0_onchip_ram_s1_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	signal mm_interconnect_0_onchip_ram_s1_write                           : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	signal mm_interconnect_0_onchip_ram_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	signal mm_interconnect_0_onchip_ram_s1_clken                           : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	signal mm_interconnect_0_descriptor_memory_s1_chipselect               : std_logic;                     -- mm_interconnect_0:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	signal mm_interconnect_0_descriptor_memory_s1_readdata                 : std_logic_vector(31 downto 0); -- descriptor_memory:readdata -> mm_interconnect_0:descriptor_memory_s1_readdata
	signal mm_interconnect_0_descriptor_memory_s1_address                  : std_logic_vector(10 downto 0); -- mm_interconnect_0:descriptor_memory_s1_address -> descriptor_memory:address
	signal mm_interconnect_0_descriptor_memory_s1_byteenable               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	signal mm_interconnect_0_descriptor_memory_s1_write                    : std_logic;                     -- mm_interconnect_0:descriptor_memory_s1_write -> descriptor_memory:write
	signal mm_interconnect_0_descriptor_memory_s1_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	signal mm_interconnect_0_descriptor_memory_s1_clken                    : std_logic;                     -- mm_interconnect_0:descriptor_memory_s1_clken -> descriptor_memory:clken
	signal mm_interconnect_0_onchip_ram_s2_chipselect                      : std_logic;                     -- mm_interconnect_0:onchip_ram_s2_chipselect -> onchip_ram:chipselect2
	signal mm_interconnect_0_onchip_ram_s2_readdata                        : std_logic_vector(31 downto 0); -- onchip_ram:readdata2 -> mm_interconnect_0:onchip_ram_s2_readdata
	signal mm_interconnect_0_onchip_ram_s2_address                         : std_logic_vector(18 downto 0); -- mm_interconnect_0:onchip_ram_s2_address -> onchip_ram:address2
	signal mm_interconnect_0_onchip_ram_s2_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_ram_s2_byteenable -> onchip_ram:byteenable2
	signal mm_interconnect_0_onchip_ram_s2_write                           : std_logic;                     -- mm_interconnect_0:onchip_ram_s2_write -> onchip_ram:write2
	signal mm_interconnect_0_onchip_ram_s2_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_ram_s2_writedata -> onchip_ram:writedata2
	signal mm_interconnect_0_onchip_ram_s2_clken                           : std_logic;                     -- mm_interconnect_0:onchip_ram_s2_clken -> onchip_ram:clken2
	signal mm_interconnect_0_ext_flash_uas_readdata                        : std_logic_vector(15 downto 0); -- ext_flash:uas_readdata -> mm_interconnect_0:ext_flash_uas_readdata
	signal mm_interconnect_0_ext_flash_uas_waitrequest                     : std_logic;                     -- ext_flash:uas_waitrequest -> mm_interconnect_0:ext_flash_uas_waitrequest
	signal mm_interconnect_0_ext_flash_uas_debugaccess                     : std_logic;                     -- mm_interconnect_0:ext_flash_uas_debugaccess -> ext_flash:uas_debugaccess
	signal mm_interconnect_0_ext_flash_uas_address                         : std_logic_vector(26 downto 0); -- mm_interconnect_0:ext_flash_uas_address -> ext_flash:uas_address
	signal mm_interconnect_0_ext_flash_uas_read                            : std_logic;                     -- mm_interconnect_0:ext_flash_uas_read -> ext_flash:uas_read
	signal mm_interconnect_0_ext_flash_uas_byteenable                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ext_flash_uas_byteenable -> ext_flash:uas_byteenable
	signal mm_interconnect_0_ext_flash_uas_readdatavalid                   : std_logic;                     -- ext_flash:uas_readdatavalid -> mm_interconnect_0:ext_flash_uas_readdatavalid
	signal mm_interconnect_0_ext_flash_uas_lock                            : std_logic;                     -- mm_interconnect_0:ext_flash_uas_lock -> ext_flash:uas_lock
	signal mm_interconnect_0_ext_flash_uas_write                           : std_logic;                     -- mm_interconnect_0:ext_flash_uas_write -> ext_flash:uas_write
	signal mm_interconnect_0_ext_flash_uas_writedata                       : std_logic_vector(15 downto 0); -- mm_interconnect_0:ext_flash_uas_writedata -> ext_flash:uas_writedata
	signal mm_interconnect_0_ext_flash_uas_burstcount                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ext_flash_uas_burstcount -> ext_flash:uas_burstcount
	signal pb_cpu_to_io_m0_waitrequest                                     : std_logic;                     -- mm_interconnect_1:pb_cpu_to_io_m0_waitrequest -> pb_cpu_to_io:m0_waitrequest
	signal pb_cpu_to_io_m0_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_1:pb_cpu_to_io_m0_readdata -> pb_cpu_to_io:m0_readdata
	signal pb_cpu_to_io_m0_debugaccess                                     : std_logic;                     -- pb_cpu_to_io:m0_debugaccess -> mm_interconnect_1:pb_cpu_to_io_m0_debugaccess
	signal pb_cpu_to_io_m0_address                                         : std_logic_vector(9 downto 0);  -- pb_cpu_to_io:m0_address -> mm_interconnect_1:pb_cpu_to_io_m0_address
	signal pb_cpu_to_io_m0_read                                            : std_logic;                     -- pb_cpu_to_io:m0_read -> mm_interconnect_1:pb_cpu_to_io_m0_read
	signal pb_cpu_to_io_m0_byteenable                                      : std_logic_vector(3 downto 0);  -- pb_cpu_to_io:m0_byteenable -> mm_interconnect_1:pb_cpu_to_io_m0_byteenable
	signal pb_cpu_to_io_m0_readdatavalid                                   : std_logic;                     -- mm_interconnect_1:pb_cpu_to_io_m0_readdatavalid -> pb_cpu_to_io:m0_readdatavalid
	signal pb_cpu_to_io_m0_writedata                                       : std_logic_vector(31 downto 0); -- pb_cpu_to_io:m0_writedata -> mm_interconnect_1:pb_cpu_to_io_m0_writedata
	signal pb_cpu_to_io_m0_write                                           : std_logic;                     -- pb_cpu_to_io:m0_write -> mm_interconnect_1:pb_cpu_to_io_m0_write
	signal pb_cpu_to_io_m0_burstcount                                      : std_logic_vector(0 downto 0);  -- pb_cpu_to_io:m0_burstcount -> mm_interconnect_1:pb_cpu_to_io_m0_burstcount
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_1_sysid_control_slave_readdata                  : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	signal mm_interconnect_1_sysid_control_slave_address                   : std_logic_vector(0 downto 0);  -- mm_interconnect_1:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_1_lcd_control_slave_readdata                    : std_logic_vector(7 downto 0);  -- lcd:readdata -> mm_interconnect_1:lcd_control_slave_readdata
	signal mm_interconnect_1_lcd_control_slave_address                     : std_logic_vector(1 downto 0);  -- mm_interconnect_1:lcd_control_slave_address -> lcd:address
	signal mm_interconnect_1_lcd_control_slave_read                        : std_logic;                     -- mm_interconnect_1:lcd_control_slave_read -> lcd:read
	signal mm_interconnect_1_lcd_control_slave_begintransfer               : std_logic;                     -- mm_interconnect_1:lcd_control_slave_begintransfer -> lcd:begintransfer
	signal mm_interconnect_1_lcd_control_slave_write                       : std_logic;                     -- mm_interconnect_1:lcd_control_slave_write -> lcd:write
	signal mm_interconnect_1_lcd_control_slave_writedata                   : std_logic_vector(7 downto 0);  -- mm_interconnect_1:lcd_control_slave_writedata -> lcd:writedata
	signal mm_interconnect_1_sys_clk_timer_s1_chipselect                   : std_logic;                     -- mm_interconnect_1:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	signal mm_interconnect_1_sys_clk_timer_s1_readdata                     : std_logic_vector(15 downto 0); -- sys_clk_timer:readdata -> mm_interconnect_1:sys_clk_timer_s1_readdata
	signal mm_interconnect_1_sys_clk_timer_s1_address                      : std_logic_vector(2 downto 0);  -- mm_interconnect_1:sys_clk_timer_s1_address -> sys_clk_timer:address
	signal mm_interconnect_1_sys_clk_timer_s1_write                        : std_logic;                     -- mm_interconnect_1:sys_clk_timer_s1_write -> mm_interconnect_1_sys_clk_timer_s1_write:in
	signal mm_interconnect_1_sys_clk_timer_s1_writedata                    : std_logic_vector(15 downto 0); -- mm_interconnect_1:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	signal mm_interconnect_1_high_res_timer_s1_chipselect                  : std_logic;                     -- mm_interconnect_1:high_res_timer_s1_chipselect -> high_res_timer:chipselect
	signal mm_interconnect_1_high_res_timer_s1_readdata                    : std_logic_vector(15 downto 0); -- high_res_timer:readdata -> mm_interconnect_1:high_res_timer_s1_readdata
	signal mm_interconnect_1_high_res_timer_s1_address                     : std_logic_vector(2 downto 0);  -- mm_interconnect_1:high_res_timer_s1_address -> high_res_timer:address
	signal mm_interconnect_1_high_res_timer_s1_write                       : std_logic;                     -- mm_interconnect_1:high_res_timer_s1_write -> mm_interconnect_1_high_res_timer_s1_write:in
	signal mm_interconnect_1_high_res_timer_s1_writedata                   : std_logic_vector(15 downto 0); -- mm_interconnect_1:high_res_timer_s1_writedata -> high_res_timer:writedata
	signal mm_interconnect_1_samplenum_s1_chipselect                       : std_logic;                     -- mm_interconnect_1:sampleNum_s1_chipselect -> sampleNum:chipselect
	signal mm_interconnect_1_samplenum_s1_readdata                         : std_logic_vector(31 downto 0); -- sampleNum:readdata -> mm_interconnect_1:sampleNum_s1_readdata
	signal mm_interconnect_1_samplenum_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_1:sampleNum_s1_address -> sampleNum:address
	signal mm_interconnect_1_samplenum_s1_write                            : std_logic;                     -- mm_interconnect_1:sampleNum_s1_write -> mm_interconnect_1_samplenum_s1_write:in
	signal mm_interconnect_1_samplenum_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_1:sampleNum_s1_writedata -> sampleNum:writedata
	signal mm_interconnect_1_adc_control_s1_chipselect                     : std_logic;                     -- mm_interconnect_1:adc_control_s1_chipselect -> adc_control:chipselect
	signal mm_interconnect_1_adc_control_s1_readdata                       : std_logic_vector(31 downto 0); -- adc_control:readdata -> mm_interconnect_1:adc_control_s1_readdata
	signal mm_interconnect_1_adc_control_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_1:adc_control_s1_address -> adc_control:address
	signal mm_interconnect_1_adc_control_s1_write                          : std_logic;                     -- mm_interconnect_1:adc_control_s1_write -> mm_interconnect_1_adc_control_s1_write:in
	signal mm_interconnect_1_adc_control_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_1:adc_control_s1_writedata -> adc_control:writedata
	signal mm_interconnect_1_wavesample_s1_readdata                        : std_logic_vector(31 downto 0); -- waveSample:readdata -> mm_interconnect_1:waveSample_s1_readdata
	signal mm_interconnect_1_wavesample_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_1:waveSample_s1_address -> waveSample:address
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- sgdma_rx:csr_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- sgdma_tx:csr_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- sys_clk_timer:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                     -- high_res_timer:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver4_irq
	signal cpu_irq_irq                                                     : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal tse_mac_receive_valid                                           : std_logic;                     -- tse_mac:ff_rx_dval -> avalon_st_adapter:in_0_valid
	signal tse_mac_receive_data                                            : std_logic_vector(31 downto 0); -- tse_mac:ff_rx_data -> avalon_st_adapter:in_0_data
	signal tse_mac_receive_ready                                           : std_logic;                     -- avalon_st_adapter:in_0_ready -> tse_mac:ff_rx_rdy
	signal tse_mac_receive_startofpacket                                   : std_logic;                     -- tse_mac:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	signal tse_mac_receive_endofpacket                                     : std_logic;                     -- tse_mac:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	signal tse_mac_receive_error                                           : std_logic_vector(5 downto 0);  -- tse_mac:rx_err -> avalon_st_adapter:in_0_error
	signal tse_mac_receive_empty                                           : std_logic_vector(1 downto 0);  -- tse_mac:ff_rx_mod -> avalon_st_adapter:in_0_empty
	signal avalon_st_adapter_out_0_valid                                   : std_logic;                     -- avalon_st_adapter:out_0_valid -> sgdma_rx:in_valid
	signal avalon_st_adapter_out_0_data                                    : std_logic_vector(31 downto 0); -- avalon_st_adapter:out_0_data -> sgdma_rx:in_data
	signal avalon_st_adapter_out_0_ready                                   : std_logic;                     -- sgdma_rx:in_ready -> avalon_st_adapter:out_0_ready
	signal avalon_st_adapter_out_0_startofpacket                           : std_logic;                     -- avalon_st_adapter:out_0_startofpacket -> sgdma_rx:in_startofpacket
	signal avalon_st_adapter_out_0_endofpacket                             : std_logic;                     -- avalon_st_adapter:out_0_endofpacket -> sgdma_rx:in_endofpacket
	signal avalon_st_adapter_out_0_error                                   : std_logic_vector(5 downto 0);  -- avalon_st_adapter:out_0_error -> sgdma_rx:in_error
	signal avalon_st_adapter_out_0_empty                                   : std_logic_vector(1 downto 0);  -- avalon_st_adapter:out_0_empty -> sgdma_rx:in_empty
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, cfi_flash_atb_bridge_0:reset, descriptor_memory:reset, ext_flash:reset_reset, mm_interconnect_0:sgdma_tx_reset_reset_bridge_in_reset_reset, mm_interconnect_1:jtag_uart_0_reset_reset_bridge_in_reset_reset, onchip_ram:reset, onchip_ram:reset2, rst_controller_reset_out_reset:in, rst_translator:in_reset, tse_mac:reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [descriptor_memory:reset_req, onchip_ram:reset_req, onchip_ram:reset_req2, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pb_cpu_to_io_reset_reset_bridge_in_reset_reset, pb_cpu_to_io:reset, rst_controller_001_reset_out_reset:in, rst_translator_001:in_reset]
	signal rst_controller_001_reset_out_reset_req                          : std_logic;                     -- rst_controller_001:reset_req -> [cpu:reset_req, rst_translator_001:reset_req_in]
	signal cpu_debug_reset_request_reset                                   : std_logic;                     -- cpu:debug_reset_request -> rst_controller_001:reset_in1
	signal merged_resets_in_reset_reset_n_ports_inv                        : std_logic;                     -- merged_resets_in_reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0, rst_controller_001:reset_in2]
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_1_sys_clk_timer_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_1_sys_clk_timer_s1_write:inv -> sys_clk_timer:write_n
	signal mm_interconnect_1_high_res_timer_s1_write_ports_inv             : std_logic;                     -- mm_interconnect_1_high_res_timer_s1_write:inv -> high_res_timer:write_n
	signal mm_interconnect_1_samplenum_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_1_samplenum_s1_write:inv -> sampleNum:write_n
	signal mm_interconnect_1_adc_control_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_1_adc_control_s1_write:inv -> adc_control:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [adc_control:reset_n, high_res_timer:reset_n, jtag_uart_0:rst_n, lcd:reset_n, sampleNum:reset_n, sgdma_rx:system_reset_n, sgdma_tx:system_reset_n, sys_clk_timer:reset_n, sysid:reset_n, waveSample:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> cpu:reset_n

begin

	adc_control : component Nios_CPU_qsys_adc_control
		port map (
			clk        => clk_clk,                                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_1_adc_control_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_adc_control_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_adc_control_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_adc_control_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_adc_control_s1_readdata,        --                    .readdata
			out_port   => adc_control_out_export                            -- external_connection.export
		);

	cfi_flash_atb_bridge_0 : component Nios_CPU_qsys_cfi_flash_atb_bridge_0
		port map (
			clk                         => clk_clk,                                         --   clk.clk
			reset                       => rst_controller_reset_out_reset,                  -- reset.reset
			request                     => ext_flash_tcm_request,                           --   tcs.request
			grant                       => ext_flash_tcm_grant,                             --      .grant
			tcs_tcm_address_out         => ext_flash_tcm_address_out,                       --      .address_out
			tcs_tcm_read_n_out(0)       => ext_flash_tcm_read_n_out,                        --      .read_n_out
			tcs_tcm_write_n_out(0)      => ext_flash_tcm_write_n_out,                       --      .write_n_out
			tcs_tcm_data_out            => ext_flash_tcm_data_out,                          --      .data_out
			tcs_tcm_data_outen          => ext_flash_tcm_data_outen,                        --      .data_outen
			tcs_tcm_data_in             => ext_flash_tcm_data_in,                           --      .data_in
			tcs_tcm_chipselect_n_out(0) => ext_flash_tcm_chipselect_n_out,                  --      .chipselect_n_out
			tcm_address_out             => cfi_flash_atb_bridge_0_out_tcm_address_out,      --   out.tcm_address_out
			tcm_read_n_out              => cfi_flash_atb_bridge_0_out_tcm_read_n_out,       --      .tcm_read_n_out
			tcm_write_n_out             => cfi_flash_atb_bridge_0_out_tcm_write_n_out,      --      .tcm_write_n_out
			tcm_data_out                => cfi_flash_atb_bridge_0_out_tcm_data_out,         --      .tcm_data_out
			tcm_chipselect_n_out        => cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out  --      .tcm_chipselect_n_out
		);

	cpu : component Nios_CPU_qsys_cpu
		port map (
			clk                                 => clk_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,      --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,            --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	descriptor_memory : component Nios_CPU_qsys_descriptor_memory
		port map (
			clk        => clk_clk,                                           --   clk1.clk
			address    => mm_interconnect_0_descriptor_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_descriptor_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_descriptor_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_descriptor_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_descriptor_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_descriptor_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_descriptor_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                    -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,                --       .reset_req
			freeze     => '0'                                                -- (terminated)
		);

	enet_pll : component Nios_CPU_qsys_enet_pll
		port map (
			refclk   => clk_clk,                --  refclk.clk
			rst      => enet_pll_reset_reset,   --   reset.reset
			outclk_0 => enet_pll_outclk0_clk,   -- outclk0.clk
			outclk_1 => enet_pll_outclk1_clk,   -- outclk1.clk
			outclk_2 => enet_pll_outclk2_clk,   -- outclk2.clk
			locked   => enet_pll_locked_export  --  locked.export
		);

	ext_flash : component Nios_CPU_qsys_ext_flash
		generic map (
			TCM_ADDRESS_W                  => 27,
			TCM_DATA_W                     => 16,
			TCM_BYTEENABLE_W               => 2,
			TCM_READ_WAIT                  => 135,
			TCM_WRITE_WAIT                 => 135,
			TCM_SETUP_WAIT                 => 25,
			TCM_DATA_HOLD                  => 20,
			TCM_TURNAROUND_TIME            => 2,
			TCM_TIMING_UNITS               => 0,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 2,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 1,
			USE_WRITE                      => 1,
			USE_BYTEENABLE                 => 0,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 0,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 0,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 0,
			ACTIVE_LOW_READ                => 1,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 1,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 0,
			ACTIVE_LOW_OUTPUTENABLE        => 0,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 1
		)
		port map (
			clk_clk              => clk_clk,                                       --   clk.clk
			reset_reset          => rst_controller_reset_out_reset,                -- reset.reset
			uas_address          => mm_interconnect_0_ext_flash_uas_address,       --   uas.address
			uas_burstcount       => mm_interconnect_0_ext_flash_uas_burstcount,    --      .burstcount
			uas_read             => mm_interconnect_0_ext_flash_uas_read,          --      .read
			uas_write            => mm_interconnect_0_ext_flash_uas_write,         --      .write
			uas_waitrequest      => mm_interconnect_0_ext_flash_uas_waitrequest,   --      .waitrequest
			uas_readdatavalid    => mm_interconnect_0_ext_flash_uas_readdatavalid, --      .readdatavalid
			uas_byteenable       => mm_interconnect_0_ext_flash_uas_byteenable,    --      .byteenable
			uas_readdata         => mm_interconnect_0_ext_flash_uas_readdata,      --      .readdata
			uas_writedata        => mm_interconnect_0_ext_flash_uas_writedata,     --      .writedata
			uas_lock             => mm_interconnect_0_ext_flash_uas_lock,          --      .lock
			uas_debugaccess      => mm_interconnect_0_ext_flash_uas_debugaccess,   --      .debugaccess
			tcm_write_n_out      => ext_flash_tcm_write_n_out,                     --   tcm.write_n_out
			tcm_read_n_out       => ext_flash_tcm_read_n_out,                      --      .read_n_out
			tcm_chipselect_n_out => ext_flash_tcm_chipselect_n_out,                --      .chipselect_n_out
			tcm_request          => ext_flash_tcm_request,                         --      .request
			tcm_grant            => ext_flash_tcm_grant,                           --      .grant
			tcm_address_out      => ext_flash_tcm_address_out,                     --      .address_out
			tcm_data_out         => ext_flash_tcm_data_out,                        --      .data_out
			tcm_data_outen       => ext_flash_tcm_data_outen,                      --      .data_outen
			tcm_data_in          => ext_flash_tcm_data_in                          --      .data_in
		);

	high_res_timer : component Nios_CPU_qsys_high_res_timer
		port map (
			clk        => clk_clk,                                             --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            -- reset.reset_n
			address    => mm_interconnect_1_high_res_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_1_high_res_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_1_high_res_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_1_high_res_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_1_high_res_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver3_irq                             --   irq.irq
		);

	jtag_uart_0 : component Nios_CPU_qsys_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver4_irq                                         --               irq.irq
		);

	lcd : component Nios_CPU_qsys_lcd
		port map (
			reset_n       => rst_controller_reset_out_reset_ports_inv,          --         reset.reset_n
			clk           => clk_clk,                                           --           clk.clk
			begintransfer => mm_interconnect_1_lcd_control_slave_begintransfer, -- control_slave.begintransfer
			read          => mm_interconnect_1_lcd_control_slave_read,          --              .read
			write         => mm_interconnect_1_lcd_control_slave_write,         --              .write
			readdata      => mm_interconnect_1_lcd_control_slave_readdata,      --              .readdata
			writedata     => mm_interconnect_1_lcd_control_slave_writedata,     --              .writedata
			address       => mm_interconnect_1_lcd_control_slave_address,       --              .address
			LCD_RS        => lcd_external_RS,                                   --      external.export
			LCD_RW        => lcd_external_RW,                                   --              .export
			LCD_data      => lcd_external_data,                                 --              .export
			LCD_E         => lcd_external_E                                     --              .export
		);

	onchip_ram : component Nios_CPU_qsys_onchip_ram
		port map (
			clk         => clk_clk,                                    --   clk1.clk
			address     => mm_interconnect_0_onchip_ram_s1_address,    --     s1.address
			clken       => mm_interconnect_0_onchip_ram_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_onchip_ram_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_onchip_ram_s1_write,      --       .write
			readdata    => mm_interconnect_0_onchip_ram_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_onchip_ram_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_onchip_ram_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,         --       .reset_req
			address2    => mm_interconnect_0_onchip_ram_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_onchip_ram_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_onchip_ram_s2_clken,      --       .clken
			write2      => mm_interconnect_0_onchip_ram_s2_write,      --       .write
			readdata2   => mm_interconnect_0_onchip_ram_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_onchip_ram_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_onchip_ram_s2_byteenable, --       .byteenable
			clk2        => clk_clk,                                    --   clk2.clk
			reset2      => rst_controller_reset_out_reset,             -- reset2.reset
			reset_req2  => rst_controller_reset_out_reset_req,         --       .reset_req
			freeze      => '0'                                         -- (terminated)
		);

	pb_cpu_to_io : component altera_avalon_mm_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 10,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => clk_clk,                                         --   clk.clk
			reset            => rst_controller_001_reset_out_reset,              -- reset.reset
			s0_waitrequest   => mm_interconnect_0_pb_cpu_to_io_s0_waitrequest,   --    s0.waitrequest
			s0_readdata      => mm_interconnect_0_pb_cpu_to_io_s0_readdata,      --      .readdata
			s0_readdatavalid => mm_interconnect_0_pb_cpu_to_io_s0_readdatavalid, --      .readdatavalid
			s0_burstcount    => mm_interconnect_0_pb_cpu_to_io_s0_burstcount,    --      .burstcount
			s0_writedata     => mm_interconnect_0_pb_cpu_to_io_s0_writedata,     --      .writedata
			s0_address       => mm_interconnect_0_pb_cpu_to_io_s0_address,       --      .address
			s0_write         => mm_interconnect_0_pb_cpu_to_io_s0_write,         --      .write
			s0_read          => mm_interconnect_0_pb_cpu_to_io_s0_read,          --      .read
			s0_byteenable    => mm_interconnect_0_pb_cpu_to_io_s0_byteenable,    --      .byteenable
			s0_debugaccess   => mm_interconnect_0_pb_cpu_to_io_s0_debugaccess,   --      .debugaccess
			m0_waitrequest   => pb_cpu_to_io_m0_waitrequest,                     --    m0.waitrequest
			m0_readdata      => pb_cpu_to_io_m0_readdata,                        --      .readdata
			m0_readdatavalid => pb_cpu_to_io_m0_readdatavalid,                   --      .readdatavalid
			m0_burstcount    => pb_cpu_to_io_m0_burstcount,                      --      .burstcount
			m0_writedata     => pb_cpu_to_io_m0_writedata,                       --      .writedata
			m0_address       => pb_cpu_to_io_m0_address,                         --      .address
			m0_write         => pb_cpu_to_io_m0_write,                           --      .write
			m0_read          => pb_cpu_to_io_m0_read,                            --      .read
			m0_byteenable    => pb_cpu_to_io_m0_byteenable,                      --      .byteenable
			m0_debugaccess   => pb_cpu_to_io_m0_debugaccess,                     --      .debugaccess
			s0_response      => open,                                            -- (terminated)
			m0_response      => "00"                                             -- (terminated)
		);

	samplenum : component Nios_CPU_qsys_sampleNum
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_1_samplenum_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_samplenum_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_samplenum_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_samplenum_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_samplenum_s1_readdata,        --                    .readdata
			out_port   => samplenum_out_export                            -- external_connection.export
		);

	sgdma_rx : component Nios_CPU_qsys_sgdma_rx
		port map (
			clk                           => clk_clk,                                   --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv,  --            reset.reset_n
			csr_chipselect                => mm_interconnect_0_sgdma_rx_csr_chipselect, --              csr.chipselect
			csr_address                   => mm_interconnect_0_sgdma_rx_csr_address,    --                 .address
			csr_read                      => mm_interconnect_0_sgdma_rx_csr_read,       --                 .read
			csr_write                     => mm_interconnect_0_sgdma_rx_csr_write,      --                 .write
			csr_writedata                 => mm_interconnect_0_sgdma_rx_csr_writedata,  --                 .writedata
			csr_readdata                  => mm_interconnect_0_sgdma_rx_csr_readdata,   --                 .readdata
			descriptor_read_readdata      => sgdma_rx_descriptor_read_readdata,         --  descriptor_read.readdata
			descriptor_read_readdatavalid => sgdma_rx_descriptor_read_readdatavalid,    --                 .readdatavalid
			descriptor_read_waitrequest   => sgdma_rx_descriptor_read_waitrequest,      --                 .waitrequest
			descriptor_read_address       => sgdma_rx_descriptor_read_address,          --                 .address
			descriptor_read_read          => sgdma_rx_descriptor_read_read,             --                 .read
			descriptor_write_waitrequest  => sgdma_rx_descriptor_write_waitrequest,     -- descriptor_write.waitrequest
			descriptor_write_address      => sgdma_rx_descriptor_write_address,         --                 .address
			descriptor_write_write        => sgdma_rx_descriptor_write_write,           --                 .write
			descriptor_write_writedata    => sgdma_rx_descriptor_write_writedata,       --                 .writedata
			csr_irq                       => irq_mapper_receiver0_irq,                  --          csr_irq.irq
			in_startofpacket              => avalon_st_adapter_out_0_startofpacket,     --               in.startofpacket
			in_endofpacket                => avalon_st_adapter_out_0_endofpacket,       --                 .endofpacket
			in_data                       => avalon_st_adapter_out_0_data,              --                 .data
			in_valid                      => avalon_st_adapter_out_0_valid,             --                 .valid
			in_ready                      => avalon_st_adapter_out_0_ready,             --                 .ready
			in_empty                      => avalon_st_adapter_out_0_empty,             --                 .empty
			in_error                      => avalon_st_adapter_out_0_error,             --                 .error
			m_write_waitrequest           => sgdma_rx_m_write_waitrequest,              --          m_write.waitrequest
			m_write_address               => sgdma_rx_m_write_address,                  --                 .address
			m_write_write                 => sgdma_rx_m_write_write,                    --                 .write
			m_write_writedata             => sgdma_rx_m_write_writedata,                --                 .writedata
			m_write_byteenable            => sgdma_rx_m_write_byteenable                --                 .byteenable
		);

	sgdma_tx : component Nios_CPU_qsys_sgdma_tx
		port map (
			clk                           => clk_clk,                                   --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv,  --            reset.reset_n
			csr_chipselect                => mm_interconnect_0_sgdma_tx_csr_chipselect, --              csr.chipselect
			csr_address                   => mm_interconnect_0_sgdma_tx_csr_address,    --                 .address
			csr_read                      => mm_interconnect_0_sgdma_tx_csr_read,       --                 .read
			csr_write                     => mm_interconnect_0_sgdma_tx_csr_write,      --                 .write
			csr_writedata                 => mm_interconnect_0_sgdma_tx_csr_writedata,  --                 .writedata
			csr_readdata                  => mm_interconnect_0_sgdma_tx_csr_readdata,   --                 .readdata
			descriptor_read_readdata      => sgdma_tx_descriptor_read_readdata,         --  descriptor_read.readdata
			descriptor_read_readdatavalid => sgdma_tx_descriptor_read_readdatavalid,    --                 .readdatavalid
			descriptor_read_waitrequest   => sgdma_tx_descriptor_read_waitrequest,      --                 .waitrequest
			descriptor_read_address       => sgdma_tx_descriptor_read_address,          --                 .address
			descriptor_read_read          => sgdma_tx_descriptor_read_read,             --                 .read
			descriptor_write_waitrequest  => sgdma_tx_descriptor_write_waitrequest,     -- descriptor_write.waitrequest
			descriptor_write_address      => sgdma_tx_descriptor_write_address,         --                 .address
			descriptor_write_write        => sgdma_tx_descriptor_write_write,           --                 .write
			descriptor_write_writedata    => sgdma_tx_descriptor_write_writedata,       --                 .writedata
			csr_irq                       => irq_mapper_receiver1_irq,                  --          csr_irq.irq
			m_read_readdata               => sgdma_tx_m_read_readdata,                  --           m_read.readdata
			m_read_readdatavalid          => sgdma_tx_m_read_readdatavalid,             --                 .readdatavalid
			m_read_waitrequest            => sgdma_tx_m_read_waitrequest,               --                 .waitrequest
			m_read_address                => sgdma_tx_m_read_address,                   --                 .address
			m_read_read                   => sgdma_tx_m_read_read,                      --                 .read
			out_data                      => sgdma_tx_out_data,                         --              out.data
			out_valid                     => sgdma_tx_out_valid,                        --                 .valid
			out_ready                     => sgdma_tx_out_ready,                        --                 .ready
			out_endofpacket               => sgdma_tx_out_endofpacket,                  --                 .endofpacket
			out_startofpacket             => sgdma_tx_out_startofpacket,                --                 .startofpacket
			out_empty                     => sgdma_tx_out_empty,                        --                 .empty
			out_error                     => sgdma_tx_out_error                         --                 .error
		);

	sys_clk_timer : component Nios_CPU_qsys_sys_clk_timer
		port map (
			clk        => clk_clk,                                            --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           -- reset.reset_n
			address    => mm_interconnect_1_sys_clk_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_1_sys_clk_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_1_sys_clk_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_1_sys_clk_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_1_sys_clk_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                            --   irq.irq
		);

	sysid : component Nios_CPU_qsys_sysid
		port map (
			clock    => clk_clk,                                          --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_1_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_1_sysid_control_slave_address(0)  --              .address
		);

	tse_mac : component Nios_CPU_qsys_tse_mac
		port map (
			clk           => clk_clk,                                            -- control_port_clock_connection.clk
			reset         => rst_controller_reset_out_reset,                     --              reset_connection.reset
			reg_addr      => mm_interconnect_0_tse_mac_control_port_address,     --                  control_port.address
			reg_data_out  => mm_interconnect_0_tse_mac_control_port_readdata,    --                              .readdata
			reg_rd        => mm_interconnect_0_tse_mac_control_port_read,        --                              .read
			reg_data_in   => mm_interconnect_0_tse_mac_control_port_writedata,   --                              .writedata
			reg_wr        => mm_interconnect_0_tse_mac_control_port_write,       --                              .write
			reg_busy      => mm_interconnect_0_tse_mac_control_port_waitrequest, --                              .waitrequest
			tx_clk        => tse_mac_pcs_mac_tx_clock_connection_clk,            --   pcs_mac_tx_clock_connection.clk
			rx_clk        => tse_mac_pcs_mac_rx_clock_connection_clk,            --   pcs_mac_rx_clock_connection.clk
			set_10        => tse_mac_mac_status_connection_set_10,               --         mac_status_connection.set_10
			set_1000      => tse_mac_mac_status_connection_set_1000,             --                              .set_1000
			eth_mode      => tse_mac_mac_status_connection_eth_mode,             --                              .eth_mode
			ena_10        => tse_mac_mac_status_connection_ena_10,               --                              .ena_10
			rgmii_in      => tse_mac_mac_rgmii_connection_rgmii_in,              --          mac_rgmii_connection.rgmii_in
			rgmii_out     => tse_mac_mac_rgmii_connection_rgmii_out,             --                              .rgmii_out
			rx_control    => tse_mac_mac_rgmii_connection_rx_control,            --                              .rx_control
			tx_control    => tse_mac_mac_rgmii_connection_tx_control,            --                              .tx_control
			ff_rx_clk     => clk_clk,                                            --      receive_clock_connection.clk
			ff_tx_clk     => clk_clk,                                            --     transmit_clock_connection.clk
			ff_rx_data    => tse_mac_receive_data,                               --                       receive.data
			ff_rx_eop     => tse_mac_receive_endofpacket,                        --                              .endofpacket
			rx_err        => tse_mac_receive_error,                              --                              .error
			ff_rx_mod     => tse_mac_receive_empty,                              --                              .empty
			ff_rx_rdy     => tse_mac_receive_ready,                              --                              .ready
			ff_rx_sop     => tse_mac_receive_startofpacket,                      --                              .startofpacket
			ff_rx_dval    => tse_mac_receive_valid,                              --                              .valid
			ff_tx_data    => sgdma_tx_out_data,                                  --                      transmit.data
			ff_tx_eop     => sgdma_tx_out_endofpacket,                           --                              .endofpacket
			ff_tx_err     => sgdma_tx_out_error,                                 --                              .error
			ff_tx_mod     => sgdma_tx_out_empty,                                 --                              .empty
			ff_tx_rdy     => sgdma_tx_out_ready,                                 --                              .ready
			ff_tx_sop     => sgdma_tx_out_startofpacket,                         --                              .startofpacket
			ff_tx_wren    => sgdma_tx_out_valid,                                 --                              .valid
			mdc           => tse_mac_mac_mdio_connection_mdc,                    --           mac_mdio_connection.mdc
			mdio_in       => tse_mac_mac_mdio_connection_mdio_in,                --                              .mdio_in
			mdio_out      => tse_mac_mac_mdio_connection_mdio_out,               --                              .mdio_out
			mdio_oen      => tse_mac_mac_mdio_connection_mdio_oen,               --                              .mdio_oen
			xon_gen       => open,                                               --           mac_misc_connection.xon_gen
			xoff_gen      => open,                                               --                              .xoff_gen
			ff_tx_crc_fwd => open,                                               --                              .ff_tx_crc_fwd
			ff_tx_septy   => open,                                               --                              .ff_tx_septy
			tx_ff_uflow   => open,                                               --                              .tx_ff_uflow
			ff_tx_a_full  => open,                                               --                              .ff_tx_a_full
			ff_tx_a_empty => open,                                               --                              .ff_tx_a_empty
			rx_err_stat   => open,                                               --                              .rx_err_stat
			rx_frm_type   => open,                                               --                              .rx_frm_type
			ff_rx_dsav    => open,                                               --                              .ff_rx_dsav
			ff_rx_a_full  => open,                                               --                              .ff_rx_a_full
			ff_rx_a_empty => open                                                --                              .ff_rx_a_empty
		);

	wavesample : component Nios_CPU_qsys_waveSample
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_1_wavesample_s1_address,  --                  s1.address
			readdata => mm_interconnect_1_wavesample_s1_readdata, --                    .readdata
			in_port  => wavesample_in_export                      -- external_connection.export
		);

	mm_interconnect_0 : component Nios_CPU_qsys_mm_interconnect_0
		port map (
			clkin_50_clk_clk                           => clk_clk,                                            --                         clkin_50_clk.clk
			cpu_reset_reset_bridge_in_reset_reset      => rst_controller_001_reset_out_reset,                 --      cpu_reset_reset_bridge_in_reset.reset
			sgdma_tx_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                     -- sgdma_tx_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                    => cpu_data_master_address,                            --                      cpu_data_master.address
			cpu_data_master_waitrequest                => cpu_data_master_waitrequest,                        --                                     .waitrequest
			cpu_data_master_byteenable                 => cpu_data_master_byteenable,                         --                                     .byteenable
			cpu_data_master_read                       => cpu_data_master_read,                               --                                     .read
			cpu_data_master_readdata                   => cpu_data_master_readdata,                           --                                     .readdata
			cpu_data_master_readdatavalid              => cpu_data_master_readdatavalid,                      --                                     .readdatavalid
			cpu_data_master_write                      => cpu_data_master_write,                              --                                     .write
			cpu_data_master_writedata                  => cpu_data_master_writedata,                          --                                     .writedata
			cpu_data_master_debugaccess                => cpu_data_master_debugaccess,                        --                                     .debugaccess
			cpu_instruction_master_address             => cpu_instruction_master_address,                     --               cpu_instruction_master.address
			cpu_instruction_master_waitrequest         => cpu_instruction_master_waitrequest,                 --                                     .waitrequest
			cpu_instruction_master_read                => cpu_instruction_master_read,                        --                                     .read
			cpu_instruction_master_readdata            => cpu_instruction_master_readdata,                    --                                     .readdata
			cpu_instruction_master_readdatavalid       => cpu_instruction_master_readdatavalid,               --                                     .readdatavalid
			sgdma_rx_descriptor_read_address           => sgdma_rx_descriptor_read_address,                   --             sgdma_rx_descriptor_read.address
			sgdma_rx_descriptor_read_waitrequest       => sgdma_rx_descriptor_read_waitrequest,               --                                     .waitrequest
			sgdma_rx_descriptor_read_read              => sgdma_rx_descriptor_read_read,                      --                                     .read
			sgdma_rx_descriptor_read_readdata          => sgdma_rx_descriptor_read_readdata,                  --                                     .readdata
			sgdma_rx_descriptor_read_readdatavalid     => sgdma_rx_descriptor_read_readdatavalid,             --                                     .readdatavalid
			sgdma_rx_descriptor_write_address          => sgdma_rx_descriptor_write_address,                  --            sgdma_rx_descriptor_write.address
			sgdma_rx_descriptor_write_waitrequest      => sgdma_rx_descriptor_write_waitrequest,              --                                     .waitrequest
			sgdma_rx_descriptor_write_write            => sgdma_rx_descriptor_write_write,                    --                                     .write
			sgdma_rx_descriptor_write_writedata        => sgdma_rx_descriptor_write_writedata,                --                                     .writedata
			sgdma_rx_m_write_address                   => sgdma_rx_m_write_address,                           --                     sgdma_rx_m_write.address
			sgdma_rx_m_write_waitrequest               => sgdma_rx_m_write_waitrequest,                       --                                     .waitrequest
			sgdma_rx_m_write_byteenable                => sgdma_rx_m_write_byteenable,                        --                                     .byteenable
			sgdma_rx_m_write_write                     => sgdma_rx_m_write_write,                             --                                     .write
			sgdma_rx_m_write_writedata                 => sgdma_rx_m_write_writedata,                         --                                     .writedata
			sgdma_tx_descriptor_read_address           => sgdma_tx_descriptor_read_address,                   --             sgdma_tx_descriptor_read.address
			sgdma_tx_descriptor_read_waitrequest       => sgdma_tx_descriptor_read_waitrequest,               --                                     .waitrequest
			sgdma_tx_descriptor_read_read              => sgdma_tx_descriptor_read_read,                      --                                     .read
			sgdma_tx_descriptor_read_readdata          => sgdma_tx_descriptor_read_readdata,                  --                                     .readdata
			sgdma_tx_descriptor_read_readdatavalid     => sgdma_tx_descriptor_read_readdatavalid,             --                                     .readdatavalid
			sgdma_tx_descriptor_write_address          => sgdma_tx_descriptor_write_address,                  --            sgdma_tx_descriptor_write.address
			sgdma_tx_descriptor_write_waitrequest      => sgdma_tx_descriptor_write_waitrequest,              --                                     .waitrequest
			sgdma_tx_descriptor_write_write            => sgdma_tx_descriptor_write_write,                    --                                     .write
			sgdma_tx_descriptor_write_writedata        => sgdma_tx_descriptor_write_writedata,                --                                     .writedata
			sgdma_tx_m_read_address                    => sgdma_tx_m_read_address,                            --                      sgdma_tx_m_read.address
			sgdma_tx_m_read_waitrequest                => sgdma_tx_m_read_waitrequest,                        --                                     .waitrequest
			sgdma_tx_m_read_read                       => sgdma_tx_m_read_read,                               --                                     .read
			sgdma_tx_m_read_readdata                   => sgdma_tx_m_read_readdata,                           --                                     .readdata
			sgdma_tx_m_read_readdatavalid              => sgdma_tx_m_read_readdatavalid,                      --                                     .readdatavalid
			cpu_debug_mem_slave_address                => mm_interconnect_0_cpu_debug_mem_slave_address,      --                  cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                  => mm_interconnect_0_cpu_debug_mem_slave_write,        --                                     .write
			cpu_debug_mem_slave_read                   => mm_interconnect_0_cpu_debug_mem_slave_read,         --                                     .read
			cpu_debug_mem_slave_readdata               => mm_interconnect_0_cpu_debug_mem_slave_readdata,     --                                     .readdata
			cpu_debug_mem_slave_writedata              => mm_interconnect_0_cpu_debug_mem_slave_writedata,    --                                     .writedata
			cpu_debug_mem_slave_byteenable             => mm_interconnect_0_cpu_debug_mem_slave_byteenable,   --                                     .byteenable
			cpu_debug_mem_slave_waitrequest            => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,  --                                     .waitrequest
			cpu_debug_mem_slave_debugaccess            => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,  --                                     .debugaccess
			descriptor_memory_s1_address               => mm_interconnect_0_descriptor_memory_s1_address,     --                 descriptor_memory_s1.address
			descriptor_memory_s1_write                 => mm_interconnect_0_descriptor_memory_s1_write,       --                                     .write
			descriptor_memory_s1_readdata              => mm_interconnect_0_descriptor_memory_s1_readdata,    --                                     .readdata
			descriptor_memory_s1_writedata             => mm_interconnect_0_descriptor_memory_s1_writedata,   --                                     .writedata
			descriptor_memory_s1_byteenable            => mm_interconnect_0_descriptor_memory_s1_byteenable,  --                                     .byteenable
			descriptor_memory_s1_chipselect            => mm_interconnect_0_descriptor_memory_s1_chipselect,  --                                     .chipselect
			descriptor_memory_s1_clken                 => mm_interconnect_0_descriptor_memory_s1_clken,       --                                     .clken
			ext_flash_uas_address                      => mm_interconnect_0_ext_flash_uas_address,            --                        ext_flash_uas.address
			ext_flash_uas_write                        => mm_interconnect_0_ext_flash_uas_write,              --                                     .write
			ext_flash_uas_read                         => mm_interconnect_0_ext_flash_uas_read,               --                                     .read
			ext_flash_uas_readdata                     => mm_interconnect_0_ext_flash_uas_readdata,           --                                     .readdata
			ext_flash_uas_writedata                    => mm_interconnect_0_ext_flash_uas_writedata,          --                                     .writedata
			ext_flash_uas_burstcount                   => mm_interconnect_0_ext_flash_uas_burstcount,         --                                     .burstcount
			ext_flash_uas_byteenable                   => mm_interconnect_0_ext_flash_uas_byteenable,         --                                     .byteenable
			ext_flash_uas_readdatavalid                => mm_interconnect_0_ext_flash_uas_readdatavalid,      --                                     .readdatavalid
			ext_flash_uas_waitrequest                  => mm_interconnect_0_ext_flash_uas_waitrequest,        --                                     .waitrequest
			ext_flash_uas_lock                         => mm_interconnect_0_ext_flash_uas_lock,               --                                     .lock
			ext_flash_uas_debugaccess                  => mm_interconnect_0_ext_flash_uas_debugaccess,        --                                     .debugaccess
			onchip_ram_s1_address                      => mm_interconnect_0_onchip_ram_s1_address,            --                        onchip_ram_s1.address
			onchip_ram_s1_write                        => mm_interconnect_0_onchip_ram_s1_write,              --                                     .write
			onchip_ram_s1_readdata                     => mm_interconnect_0_onchip_ram_s1_readdata,           --                                     .readdata
			onchip_ram_s1_writedata                    => mm_interconnect_0_onchip_ram_s1_writedata,          --                                     .writedata
			onchip_ram_s1_byteenable                   => mm_interconnect_0_onchip_ram_s1_byteenable,         --                                     .byteenable
			onchip_ram_s1_chipselect                   => mm_interconnect_0_onchip_ram_s1_chipselect,         --                                     .chipselect
			onchip_ram_s1_clken                        => mm_interconnect_0_onchip_ram_s1_clken,              --                                     .clken
			onchip_ram_s2_address                      => mm_interconnect_0_onchip_ram_s2_address,            --                        onchip_ram_s2.address
			onchip_ram_s2_write                        => mm_interconnect_0_onchip_ram_s2_write,              --                                     .write
			onchip_ram_s2_readdata                     => mm_interconnect_0_onchip_ram_s2_readdata,           --                                     .readdata
			onchip_ram_s2_writedata                    => mm_interconnect_0_onchip_ram_s2_writedata,          --                                     .writedata
			onchip_ram_s2_byteenable                   => mm_interconnect_0_onchip_ram_s2_byteenable,         --                                     .byteenable
			onchip_ram_s2_chipselect                   => mm_interconnect_0_onchip_ram_s2_chipselect,         --                                     .chipselect
			onchip_ram_s2_clken                        => mm_interconnect_0_onchip_ram_s2_clken,              --                                     .clken
			pb_cpu_to_io_s0_address                    => mm_interconnect_0_pb_cpu_to_io_s0_address,          --                      pb_cpu_to_io_s0.address
			pb_cpu_to_io_s0_write                      => mm_interconnect_0_pb_cpu_to_io_s0_write,            --                                     .write
			pb_cpu_to_io_s0_read                       => mm_interconnect_0_pb_cpu_to_io_s0_read,             --                                     .read
			pb_cpu_to_io_s0_readdata                   => mm_interconnect_0_pb_cpu_to_io_s0_readdata,         --                                     .readdata
			pb_cpu_to_io_s0_writedata                  => mm_interconnect_0_pb_cpu_to_io_s0_writedata,        --                                     .writedata
			pb_cpu_to_io_s0_burstcount                 => mm_interconnect_0_pb_cpu_to_io_s0_burstcount,       --                                     .burstcount
			pb_cpu_to_io_s0_byteenable                 => mm_interconnect_0_pb_cpu_to_io_s0_byteenable,       --                                     .byteenable
			pb_cpu_to_io_s0_readdatavalid              => mm_interconnect_0_pb_cpu_to_io_s0_readdatavalid,    --                                     .readdatavalid
			pb_cpu_to_io_s0_waitrequest                => mm_interconnect_0_pb_cpu_to_io_s0_waitrequest,      --                                     .waitrequest
			pb_cpu_to_io_s0_debugaccess                => mm_interconnect_0_pb_cpu_to_io_s0_debugaccess,      --                                     .debugaccess
			sgdma_rx_csr_address                       => mm_interconnect_0_sgdma_rx_csr_address,             --                         sgdma_rx_csr.address
			sgdma_rx_csr_write                         => mm_interconnect_0_sgdma_rx_csr_write,               --                                     .write
			sgdma_rx_csr_read                          => mm_interconnect_0_sgdma_rx_csr_read,                --                                     .read
			sgdma_rx_csr_readdata                      => mm_interconnect_0_sgdma_rx_csr_readdata,            --                                     .readdata
			sgdma_rx_csr_writedata                     => mm_interconnect_0_sgdma_rx_csr_writedata,           --                                     .writedata
			sgdma_rx_csr_chipselect                    => mm_interconnect_0_sgdma_rx_csr_chipselect,          --                                     .chipselect
			sgdma_tx_csr_address                       => mm_interconnect_0_sgdma_tx_csr_address,             --                         sgdma_tx_csr.address
			sgdma_tx_csr_write                         => mm_interconnect_0_sgdma_tx_csr_write,               --                                     .write
			sgdma_tx_csr_read                          => mm_interconnect_0_sgdma_tx_csr_read,                --                                     .read
			sgdma_tx_csr_readdata                      => mm_interconnect_0_sgdma_tx_csr_readdata,            --                                     .readdata
			sgdma_tx_csr_writedata                     => mm_interconnect_0_sgdma_tx_csr_writedata,           --                                     .writedata
			sgdma_tx_csr_chipselect                    => mm_interconnect_0_sgdma_tx_csr_chipselect,          --                                     .chipselect
			tse_mac_control_port_address               => mm_interconnect_0_tse_mac_control_port_address,     --                 tse_mac_control_port.address
			tse_mac_control_port_write                 => mm_interconnect_0_tse_mac_control_port_write,       --                                     .write
			tse_mac_control_port_read                  => mm_interconnect_0_tse_mac_control_port_read,        --                                     .read
			tse_mac_control_port_readdata              => mm_interconnect_0_tse_mac_control_port_readdata,    --                                     .readdata
			tse_mac_control_port_writedata             => mm_interconnect_0_tse_mac_control_port_writedata,   --                                     .writedata
			tse_mac_control_port_waitrequest           => mm_interconnect_0_tse_mac_control_port_waitrequest  --                                     .waitrequest
		);

	mm_interconnect_1 : component Nios_CPU_qsys_mm_interconnect_1
		port map (
			clkin_50_clk_clk                               => clk_clk,                                                     --                             clkin_50_clk.clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                              --  jtag_uart_0_reset_reset_bridge_in_reset.reset
			pb_cpu_to_io_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                          -- pb_cpu_to_io_reset_reset_bridge_in_reset.reset
			pb_cpu_to_io_m0_address                        => pb_cpu_to_io_m0_address,                                     --                          pb_cpu_to_io_m0.address
			pb_cpu_to_io_m0_waitrequest                    => pb_cpu_to_io_m0_waitrequest,                                 --                                         .waitrequest
			pb_cpu_to_io_m0_burstcount                     => pb_cpu_to_io_m0_burstcount,                                  --                                         .burstcount
			pb_cpu_to_io_m0_byteenable                     => pb_cpu_to_io_m0_byteenable,                                  --                                         .byteenable
			pb_cpu_to_io_m0_read                           => pb_cpu_to_io_m0_read,                                        --                                         .read
			pb_cpu_to_io_m0_readdata                       => pb_cpu_to_io_m0_readdata,                                    --                                         .readdata
			pb_cpu_to_io_m0_readdatavalid                  => pb_cpu_to_io_m0_readdatavalid,                               --                                         .readdatavalid
			pb_cpu_to_io_m0_write                          => pb_cpu_to_io_m0_write,                                       --                                         .write
			pb_cpu_to_io_m0_writedata                      => pb_cpu_to_io_m0_writedata,                                   --                                         .writedata
			pb_cpu_to_io_m0_debugaccess                    => pb_cpu_to_io_m0_debugaccess,                                 --                                         .debugaccess
			adc_control_s1_address                         => mm_interconnect_1_adc_control_s1_address,                    --                           adc_control_s1.address
			adc_control_s1_write                           => mm_interconnect_1_adc_control_s1_write,                      --                                         .write
			adc_control_s1_readdata                        => mm_interconnect_1_adc_control_s1_readdata,                   --                                         .readdata
			adc_control_s1_writedata                       => mm_interconnect_1_adc_control_s1_writedata,                  --                                         .writedata
			adc_control_s1_chipselect                      => mm_interconnect_1_adc_control_s1_chipselect,                 --                                         .chipselect
			high_res_timer_s1_address                      => mm_interconnect_1_high_res_timer_s1_address,                 --                        high_res_timer_s1.address
			high_res_timer_s1_write                        => mm_interconnect_1_high_res_timer_s1_write,                   --                                         .write
			high_res_timer_s1_readdata                     => mm_interconnect_1_high_res_timer_s1_readdata,                --                                         .readdata
			high_res_timer_s1_writedata                    => mm_interconnect_1_high_res_timer_s1_writedata,               --                                         .writedata
			high_res_timer_s1_chipselect                   => mm_interconnect_1_high_res_timer_s1_chipselect,              --                                         .chipselect
			jtag_uart_0_avalon_jtag_slave_address          => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address,     --            jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write            => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write,       --                                         .write
			jtag_uart_0_avalon_jtag_slave_read             => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read,        --                                         .read
			jtag_uart_0_avalon_jtag_slave_readdata         => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata,    --                                         .readdata
			jtag_uart_0_avalon_jtag_slave_writedata        => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata,   --                                         .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest      => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                         .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect       => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                         .chipselect
			lcd_control_slave_address                      => mm_interconnect_1_lcd_control_slave_address,                 --                        lcd_control_slave.address
			lcd_control_slave_write                        => mm_interconnect_1_lcd_control_slave_write,                   --                                         .write
			lcd_control_slave_read                         => mm_interconnect_1_lcd_control_slave_read,                    --                                         .read
			lcd_control_slave_readdata                     => mm_interconnect_1_lcd_control_slave_readdata,                --                                         .readdata
			lcd_control_slave_writedata                    => mm_interconnect_1_lcd_control_slave_writedata,               --                                         .writedata
			lcd_control_slave_begintransfer                => mm_interconnect_1_lcd_control_slave_begintransfer,           --                                         .begintransfer
			sampleNum_s1_address                           => mm_interconnect_1_samplenum_s1_address,                      --                             sampleNum_s1.address
			sampleNum_s1_write                             => mm_interconnect_1_samplenum_s1_write,                        --                                         .write
			sampleNum_s1_readdata                          => mm_interconnect_1_samplenum_s1_readdata,                     --                                         .readdata
			sampleNum_s1_writedata                         => mm_interconnect_1_samplenum_s1_writedata,                    --                                         .writedata
			sampleNum_s1_chipselect                        => mm_interconnect_1_samplenum_s1_chipselect,                   --                                         .chipselect
			sys_clk_timer_s1_address                       => mm_interconnect_1_sys_clk_timer_s1_address,                  --                         sys_clk_timer_s1.address
			sys_clk_timer_s1_write                         => mm_interconnect_1_sys_clk_timer_s1_write,                    --                                         .write
			sys_clk_timer_s1_readdata                      => mm_interconnect_1_sys_clk_timer_s1_readdata,                 --                                         .readdata
			sys_clk_timer_s1_writedata                     => mm_interconnect_1_sys_clk_timer_s1_writedata,                --                                         .writedata
			sys_clk_timer_s1_chipselect                    => mm_interconnect_1_sys_clk_timer_s1_chipselect,               --                                         .chipselect
			sysid_control_slave_address                    => mm_interconnect_1_sysid_control_slave_address,               --                      sysid_control_slave.address
			sysid_control_slave_readdata                   => mm_interconnect_1_sysid_control_slave_readdata,              --                                         .readdata
			waveSample_s1_address                          => mm_interconnect_1_wavesample_s1_address,                     --                            waveSample_s1.address
			waveSample_s1_readdata                         => mm_interconnect_1_wavesample_s1_readdata                     --                                         .readdata
		);

	irq_mapper : component Nios_CPU_qsys_irq_mapper
		port map (
			clk           => clk_clk,                            --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			sender_irq    => cpu_irq_irq                         --    sender.irq
		);

	avalon_st_adapter : component Nios_CPU_qsys_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 6,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 2,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 6,
			outUseEmptyPort => 1,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => clk_clk,                               -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,        -- in_rst_0.reset
			in_0_data           => tse_mac_receive_data,                  --     in_0.data
			in_0_valid          => tse_mac_receive_valid,                 --         .valid
			in_0_ready          => tse_mac_receive_ready,                 --         .ready
			in_0_startofpacket  => tse_mac_receive_startofpacket,         --         .startofpacket
			in_0_endofpacket    => tse_mac_receive_endofpacket,           --         .endofpacket
			in_0_empty          => tse_mac_receive_empty,                 --         .empty
			in_0_error          => tse_mac_receive_error,                 --         .error
			out_0_data          => avalon_st_adapter_out_0_data,          --    out_0.data
			out_0_valid         => avalon_st_adapter_out_0_valid,         --         .valid
			out_0_ready         => avalon_st_adapter_out_0_ready,         --         .ready
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket,   --         .endofpacket
			out_0_empty         => avalon_st_adapter_out_0_empty,         --         .empty
			out_0_error         => avalon_st_adapter_out_0_error          --         .error
		);

	rst_controller : component nios_cpu_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => merged_resets_in_reset_reset_n_ports_inv, -- reset_in0.reset
			reset_in1      => merged_resets_in_reset_reset_n_ports_inv, -- reset_in1.reset
			clk            => clk_clk,                                  --       clk.clk
			reset_out      => rst_controller_reset_out_reset,           -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,       --          .reset_req
			reset_req_in0  => '0',                                      -- (terminated)
			reset_req_in1  => '0',                                      -- (terminated)
			reset_in2      => '0',                                      -- (terminated)
			reset_req_in2  => '0',                                      -- (terminated)
			reset_in3      => '0',                                      -- (terminated)
			reset_req_in3  => '0',                                      -- (terminated)
			reset_in4      => '0',                                      -- (terminated)
			reset_req_in4  => '0',                                      -- (terminated)
			reset_in5      => '0',                                      -- (terminated)
			reset_req_in5  => '0',                                      -- (terminated)
			reset_in6      => '0',                                      -- (terminated)
			reset_req_in6  => '0',                                      -- (terminated)
			reset_in7      => '0',                                      -- (terminated)
			reset_req_in7  => '0',                                      -- (terminated)
			reset_in8      => '0',                                      -- (terminated)
			reset_req_in8  => '0',                                      -- (terminated)
			reset_in9      => '0',                                      -- (terminated)
			reset_req_in9  => '0',                                      -- (terminated)
			reset_in10     => '0',                                      -- (terminated)
			reset_req_in10 => '0',                                      -- (terminated)
			reset_in11     => '0',                                      -- (terminated)
			reset_req_in11 => '0',                                      -- (terminated)
			reset_in12     => '0',                                      -- (terminated)
			reset_req_in12 => '0',                                      -- (terminated)
			reset_in13     => '0',                                      -- (terminated)
			reset_req_in13 => '0',                                      -- (terminated)
			reset_in14     => '0',                                      -- (terminated)
			reset_req_in14 => '0',                                      -- (terminated)
			reset_in15     => '0',                                      -- (terminated)
			reset_req_in15 => '0'                                       -- (terminated)
		);

	rst_controller_001 : component nios_cpu_qsys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => merged_resets_in_reset_reset_n_ports_inv, -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,            -- reset_in1.reset
			reset_in2      => merged_resets_in_reset_reset_n_ports_inv, -- reset_in2.reset
			clk            => clk_clk,                                  --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,       -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req,   --          .reset_req
			reset_req_in0  => '0',                                      -- (terminated)
			reset_req_in1  => '0',                                      -- (terminated)
			reset_req_in2  => '0',                                      -- (terminated)
			reset_in3      => '0',                                      -- (terminated)
			reset_req_in3  => '0',                                      -- (terminated)
			reset_in4      => '0',                                      -- (terminated)
			reset_req_in4  => '0',                                      -- (terminated)
			reset_in5      => '0',                                      -- (terminated)
			reset_req_in5  => '0',                                      -- (terminated)
			reset_in6      => '0',                                      -- (terminated)
			reset_req_in6  => '0',                                      -- (terminated)
			reset_in7      => '0',                                      -- (terminated)
			reset_req_in7  => '0',                                      -- (terminated)
			reset_in8      => '0',                                      -- (terminated)
			reset_req_in8  => '0',                                      -- (terminated)
			reset_in9      => '0',                                      -- (terminated)
			reset_req_in9  => '0',                                      -- (terminated)
			reset_in10     => '0',                                      -- (terminated)
			reset_req_in10 => '0',                                      -- (terminated)
			reset_in11     => '0',                                      -- (terminated)
			reset_req_in11 => '0',                                      -- (terminated)
			reset_in12     => '0',                                      -- (terminated)
			reset_req_in12 => '0',                                      -- (terminated)
			reset_in13     => '0',                                      -- (terminated)
			reset_req_in13 => '0',                                      -- (terminated)
			reset_in14     => '0',                                      -- (terminated)
			reset_req_in14 => '0',                                      -- (terminated)
			reset_in15     => '0',                                      -- (terminated)
			reset_req_in15 => '0'                                       -- (terminated)
		);

	merged_resets_in_reset_reset_n_ports_inv <= not merged_resets_in_reset_reset_n;

	mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_1_sys_clk_timer_s1_write_ports_inv <= not mm_interconnect_1_sys_clk_timer_s1_write;

	mm_interconnect_1_high_res_timer_s1_write_ports_inv <= not mm_interconnect_1_high_res_timer_s1_write;

	mm_interconnect_1_samplenum_s1_write_ports_inv <= not mm_interconnect_1_samplenum_s1_write;

	mm_interconnect_1_adc_control_s1_write_ports_inv <= not mm_interconnect_1_adc_control_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of Nios_CPU_qsys
