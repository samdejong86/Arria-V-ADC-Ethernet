// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
bkVGBcFmDjxELOla8c7sbn/HDQEfVD5MY+ilScIEx0RmBnDNEL276Rkw4BSKyQtQ
j4S0tZ/yROo+FiPXGxXkMyEZmbILsTmC23EzXGsyrO3lgIrTSrEWfoebgQ0Xp2kI
Dus0jzdzHtvRqn3J/AbXdYagBOx7FoHbbxm6MUTlNMFTUfDBwpmYhw==
//pragma protect end_key_block
//pragma protect digest_block
9w6AebajkVXuqvVfsAHhuah1av0=
//pragma protect end_digest_block
//pragma protect data_block
TrEeKlkyyG7hsCxoxCN2tjLg6KYV85t7nMiVsgf8+J6CikKSspT8dJoQrgdsPaHj
tIbpCDEWb/LM8ZhBWlKg52yVvNnl5Kh2ug/J+yPpUVA74z/jbU7zSepiM1VDCG40
8taRCmiGENiCcF8mznpSVa+dZOene94J4wYVM8Y02lsoo5UxwEOm7d0s0/RRiJsU
5QQtSyg+i+AJmKWNh0AxiZqbGKzN1ODqSBag/iyXNAwpFeCID6CRtWPidvwGSr2P
8VZE/3NZXAq/YFy4k6vpm2HHGIYzce7TEKLc1VgqaEeWpp4ykkUJQm27iuO2h+fZ
KnkZYo1KljXpQFKXUmETpwGnVMEsFfFBNiBac0njkiyhd1JxLtmt1f4AkPaLOGcI
tCLhCO9Idl3HJVcqvbffSIZxVIUwnBJniWfr7P036f0ppacG57xENf/qeq+p6PSF
bw4SDxikOto1RL2dNwKPqp8RkM0YLT0Jcqmh69xhrq93hXYwk/s3ndGBgVr6xpnr
uN04vnAvHTYS6VRj5QILOXc3LEtoU08OMwvFTMqXl4YDo5t51OgWTnTM5S35eg9q
AkSh1JqaOLU6WSVo0DLsp2WBU7DmPKi0wUcIGmhz76j5T3of3LwrabyV5UcWFddI
8HZlH3Iek7+JUUTx8EkRb2/UO5CGoJPN2YukldvLTRIjZgUw2Q2OjaeW4Uvrq24X
mbbAJ9qy7jTCwZ+PthkPNFmY8Zt9D3CK7BHOcqEP6kfINB0P6JtGeeKMVii9Z9WU
/PiwU0lCfVnCONSETlaOVLEtWdb03yR0PEs89+Q9m2btJH9+jWAILfRUHb3L0vYf
77BkueGIlKbFBNDG2fTmSN1Qd+POEJpz0JjuHt4s1uZYb0uftqkSfw/yCV6PM+j9
5dOxLr/aul2o1X7ZVWspfuN6VHR1EzvQ8Ylnl+CnPJbdN6rwJjeXFGDx2UBgvGkD
0ZwhozWHPW/k41S8ZwHdaJjy73x9/O7S/RBil3o6TKlMJFheXVlWKyRIRmCfNcVO
St2b2w6gvivOWxNJrGnW1w4b22KBgy/jDG5Yokn7HqvH5UDjeg626zaEsPv4Y/sq
wAFlfAk0TaiphWQSEI8o8e2cqVgBV/VH72yoJLstRXWOgpTtE0eLWN9FmTHt+8hs
RG/+9iGKdyKNbOuDvsOMpdy/wOLiVbJ41C9zW18SmXX6swFDMdxY2HLvDg9pYLFm
NxHqjtEZH1w+d4HG+s84biIX/YkWSMzVMdRoWGBju/ch86GBiNYeYBnDYTC7s63H
Kf47H3HaXJpCdexITwnTLgdTXEYd8OOUmwPMnvVmQKkONvQXLj3fLti8UsbH2bK/
6nbBO916w+W2VHHdiXvHI4aKmh04VgTm0ENMNE4rqq6y1t/Y70jqzKms+L4365MT
v3mkpQu1PcQvDk1o4CmIBWuAWrh7tX98ytPiFnAgV7quR7Aaggi1uv+e9T5xig5R
foJstveAsHxA3LTME0HE1YfI3Vf+HNiFQ01KIs+nZR9kFvKp0iWCb1LkfiiWJ+Pw
e1TDR9dKZC9cXpGJFmp0PXd9Ii6OHfE4xqmw5Vwepf2UjarXlE0BImikQtwY85o/
uoCwF5qykMf04tr4TzImwH0Cxt956DELJRVdU9ZgoX5v+xF1HW0LSK/Ml7IONuDz
WbKhhev4RlpJwVcsjK6PXF+niFhLisVb48oOJyQdm/ao2UFxKzWUT6XtuR1HuIkA
HCSdJ7y85kwD5MtNYFRI77tvA9JdSqcPWU8DMdVBYWELhH0be6jBlVvCgMz4eucO
UbsREHbah/gwFgOeLkIX/jsuSk4eQcPLlWki7dWYaC7makp6qiU5TWN24kxVnm/W
56a4sXekroVYwKLZ07PnhGW8/A0neHQK/pyP+mNVqURhf7qW9ubCDLCl1SmFMCNA
pKeW8PZc1lvmgsJv9JHv6jGTKjJiPt3l4o156G5l3FHKTM+syyCUrDJDy7SWUwj3
RaYOjaxKfPXHzWkQC8mPibG0AoB95GGcP6DQgtrEK9Z/jO4kHXNt+YGA1QdKHyhT
7B0J23uDsTwIesI3Z4bXIi0i52AONFvmkwlFfYrBhHtydHKSaIp8ZxdW7Kfzjr4v
sxx8YluWdYSgzo17hJMUNpmdPK36tzWqJXkZyEAvK8Icj5hL7FCSxEhIK70K2m0/
OcFziy8nY/laRbqG5nj0U0GFKBrn/PzaIk2t4HWfZSzijLlgsFa6L8u4mHNZmrTf
evbfOOo0bdUMa3kp2LYLqYF8EW2wvwjfXfCC9skNvJ49avsMDa1qdAFy1dcFpoSQ
3yF2WsJ4utzgLOo2Z7qdEwfRDR6C9Zc10DkP+xD8UvhS91WTCsGK1MRqgjs2wyg5
7xQGEEws+1LnKxBzwsZfsmC5DpTV3YKU8xAQCCUDLyYFy+LYf2G2eAKf+wzjqMRJ
ryFIzw9/DvlARVjMmOKDqaTyjNGpNSJMJsMFDSesnuPDZO0z5dcKiQSmNlRBCV36
VqdPPlBBREE2BzWJn923B11i/I0jkGPqGILNaYTLd4j5EUwyFtD9cy4HaX3vz2Mw
qS0YB6BCRh+9G8nnrmo98jyLOgrZ/6/f83aFjPtWJKEj4iMjw6mP2fMuALOaJIWM
mFEXNwEroCSVGBjrgN1EWJrQ1pZ9jduY3vgXHywj5Ij/HbGYaRLif/YNaDkCmC8g
mqhVJPJZaykxsMvXrTYeEiZbE9JR2ps9ZmiNKtA08Q3jsAI7dLzNpZUK8XEJropi
+e/SS4GNq8beaUqOlRG8H/RqWOLg0kbgee/yN5lBPhe1EeZtltvD8wnEpIjRa0XA
IokHvE2RBRUFHiYI0hMNKTQfM+DTi71VR47/ucAACClTFeMtbMh2g/0tv36ngEJg
ljQMXA5XZ7tJjr85qL2o8YVSYhqmuIwXIC6JpBdUqFBdfSqkKX27pntS/9OU9nJn
PPF2VSij3DUqTttL8g/3RnuBUOlBsT/zw2b6HcvuB2LB2XiARD6N/qFQjjTTs2ft
VdF/1oXyRao6Qs+61kM+6M5adukyYSMCkE6buEO3rtGXCFQprc4WztiH6zOHsRcU
9CuuYvIShTFhAGls0bzKPXqCEuJlki8fbIdsrKyLkb1MQ32yyA2NfYXOPP28nh3z
Zn0+qYAUTMHrkqZsrsyCKDascQyPl1h98uEDWnSp++y+phb6ZvlITsorV4MBQYnx
TI/ia/85/Kgzo+rFGjvnZKLM0deR0ezYMLWLvVraCrIfEd+0FmaNu7Mw5z617238
EDPPthl+wv0XhafdHSAdbEx2NoXImboFAaoSeZJ6SCML8RICTYBqEi9kmFlEDSo8
VaCV5ixxcNAP43uJ4UVCqxWTrw8tMYdYHCrZR+QXqZ2yeuw6h8RFMbTxeJ2ia2Vv
N8s5NcFez0mTe3wihZTjtFzj5xEgaIP/7WwYFtwee5amTnZl/1CPutTnX4muJTgD
N7R1vpQgS48ATWKQfKU9RvI0Eim3txguHowcdJqwwUvdumqD9Z3i4610bjjzTTdj
Jw8DUiGIFkFEOzL5WXpFc5m023oT8lCXG6gCT+XzAhRvjsUxpO9SGKv2jRZXh76u
K2Yh9RDJtWvAKJSHzXFr7LqaHR3ZQOlW0fJUf4sUtk8ixKWqWN0rAT2Aipp7Iqiy
kGs4e33HQi/JMns0j/B5B8CiYzm9d5tDbe2zUsH7YLjrkD2CzdbxvxKDEiR1P/cW
uLrtym8D9vu54TtCn7g6ah+yjuxe2U2NHCgDCZwfmfjxd7oZujiZiZHFcGBwC8S4
ghMpS4IeLNW5SQ7sQ1zaGwog+xZc7PUXMi4o6KQVd/FLWVP6hpPKPE+jEcF7AzZ5
QT++pOQC+kYRPUbXPCcc6YT1h6PfMFXIoRlpCKxoLNCVfVS+U7w8oOQhOMDyDL8B
ZyJ2DaQRfWuAbx4eS9sg6OjyXUGSyL64s3jr22HELt8QHBy20Kk0Tm/W8elDOLV4
unvOlpELtNWukc7K98DHGnE87L87eITZ8wIqtRS3Mw10DQeOBL0dr1Oh2Rf+GkJg
Q44DWI/ZPO1d5A6AIMJPSOku9QSNWfVgeb5/SEDLGXFOaWM7KBRIXxPJZwfzMtU/
8OZze1dhhZjJioaF5uPrk7BfGo2D/JyIn/lDwWKVD148rCL/t16xFXU+LE0ztreC
JN51rAgEHQ9NnsK3qDyQutZxuOUONIdHmepv8CmKATbs3TMbZg8zKc7FswMta74U
0QClXPf4QRfTVvKF00cH+Hju5TZRecrIbzIFiRp8TDPd8rWZuwukN+RtbG/kfqoD
StvJysMjzV2MYSMedGP6XiRV/z892r4JpbBrP1zdWK9hsbR48gmf02AHd5wtVb2t
YhBzKnU3nIXr/AnboWRYdHoZP4OWIFb7XO1jqiVSxxR8MAjIZpxjyM6EQsB4roEW
pZdgQwklbxRTqET8IHayLa3px8hz9Ny5XdaVEaClrPtoU6OjkiFbaJKYBfYjivyz
r97xeTFfNZDUNxVZEXNB+y3IaEHHJjBgPq081hgftgyDMf7218bUuZfWqMt3tRxs
ZS6VRnwdbTYxSroWThFnM3TxJyOE/TZ+6wCIqpsY4tpGgu8d3WfxFV7zGmct2kLz
kkaZ6ngwXowq2LPrOnIpHelAOdrb9vLh88P7rLXOsx2oOlmkIgXZDmXIqMmdfSQ9
20Lb39GLcgl4t37q4qu15+YfD9Diqr9Me0vuJnXAzxHu1Lb8YkxMGbZPBOCso5cW
khcYm0/7utJscFoBI9lH6lmZfrTg2OXE5dra80aCtd52m4RGpfx5wVIkYnQILuX+
zAibZVawo1YcMA3W0e2OU2PY1chKjAiTIyT9xaPfyq/9O943WdHnnZUXMrplzoEf
USHhCOglUpWXpLGtUE9e0TKwHoAqej5eKH8tzJYocBhLuBDG6fGZCrEZhABLR/kP
0pWo/K0ePUwQRV7f4g+NEWi/l5jmAvrZqB8M1qgjkSaX5taBe5PaZmCoYf4ctk3e
nPaISgQjsHtgygjFfcr7+ym2lFpkF2PcPXfTalnsrUpcsaB8dwfooth3z89DReq6
RjXxfwzSTfjeC8P9NnY58yVNyThQ2t+at9Fryvh7c0BHaHhAcYIRMo7coXwjL6Kb
8tSUjSbihdBNUutnOOJJfXfcwNPYpzGE8kJLMqpjl8MSo1eXy5eFihUpaZvyvuJ4
C0Hd7UoN3KBBBzrFLMIxPcBEceXJ0LELbroQJtQ4yWgdFmpRD3sE2CEiK3KwwKFF
oYAV4I8mhAiXbHE1kjN6Oez1PDy00eEf/kzchtN+8WHIKJjNoLf5hYTYr4HbUUqH
Rf9CGtqjNyqX+KcNaNYgZwxIdTrhoK1J4Htsx4Y5+qUc2YpUtAmxXPo8NkpYOd+W
jqlvvGbUCMgUTM96StTyoS7s0+SOdTAO+CFXgPZR1byG4uEPGAM/UCQW2sYKkGGn
zpec+sBP7rfG+aBW8Uzdeemk1f009s09y0ODHejIXZJoTCJQgu4D+6lddekoOgmA
TvxYKBXvCUKkpojTyp1Zf0YtbI00FlZTsDNpa5h2U6k6wYfoIntU+VzwaugEgX/b
31u1B1bixb9TzNHJIQ0mpmAyI/+2YTg36yFnNCJACa0iXulRYWpkRwYTuXed7H4f
MLvSHCCAqYw4LOfUWkzX0Dtw62W9OLqhwsrjA9H/h7eSEzsb2VQWwd4BUKFtoOA5
yZrEyaBQcMuOoKY4QcFkMFfZTODtnLzu4Fd3CYrMo28Gvhe40CFbcwuKxe3Aw6BQ
3+ieFOSzppl249ixBouqBB2A1t2AylxR0dDXWlKnrzhSbg0RXXaf5Qhpe3jj14+F
9gqAzYKzXfBkTe7iA74UfPonTFaAdxCJHOrrSwWdDDh7S5XezRECiWTU9LEax4Io
yrq/ydWaQaz4WvjLK68S9DSiasfk1Rwx4Ny2V9t/KfOMvja1W1vgaoqeOFQMPgr+
ruT01/HoM5GGWINANAEfiRiiv5dGiFbSHAr/cGw+CvLM+ytv78zVY0BJz+lRF/pt
9Dyxiv0ad9PE2JxsHJFmZK4PKESbTI1C3PP8x0aaJovjgu+i8XwSz1aV1cXQ4+Ct
i4EoAuA9vYpWCd3H1n0xs0Xsh69+sCd8H8hsLm0aSLvu+SHhGOqwTkWUZaohVxZa
RqWM/ZjHH2Fd7Nug41P+G7Ki9mwapLfxqNikFu9QoUKjjVJqPJwd5X6kBeszU8Y7
qFzPS/R9RJEJAGVffPZejTythVvLyZG3Cll6fXoQH5Ej9bO6SEKLRJdTdgUujXvR
wX8bkPf+wyQ0Fcyu9CCECRxhsR16lhzl2vT44+9Cz4GD1930laVU0DdaJOZoJlkN
QOwmzwVFZU4sq2gqt/LzgmYafSPXqL3Dc/nWggaPAwsTO3CSjG7tNPJjVx4gJ37f
TR6LRsrDSgu2VP7GIglU6FdHBiZmQxgzOiIEIFlMb61z8M6nF6s2VrubVedZXBmc
aYFhwjZWPdJduoTvoL7i/qiTJh+mfZ6hGJZG4UP8oTh59I6EekLBF7/c/T4znayk
mZxcj4ZG0OXmq6vcLsGYlNs57Ged8fdO7329HLpX2CgTchphJiqtLhADHjetO9k8
NuzdhM0yNp1+v0JAEjymVYcjH4tZHl78JtV+sVFNZYP0cO+UebaWPlIQ3nhsn9TZ
/x8LXd7NDL1jlPE1fFvXgDuuxvIQK+av6O8bor9rK8kGkn38Asi+yU62EQ+FjV1w
pPZ89hTU4r7VdwqPX5qQsqHcSrBLyGU59wqBvaEMg63ua9idEoIZMqctdnplnXPh
Pxr9/jTatxkfS06hWjgMegtfeSv0v8sARl5UDhIZCPXbwM2GnVmrASyDZN6i1URI
X7l7RvB18ksFay/9y+Yu3wTVyIOtBZlrPbqVlbiYJXqvgSfEguRj3vY4g8hbScY7
4dv2YQwIzcITgkVaOCucwS22TmLXqQvxT9S2dVULQhEZQqCvPPh6l5CqWD7zvqei
y9kWUn5/cUIxd/Ird09vDPtP2Wcv6UZ31NKpkAIrv34DbYie2vTvlVB1dlMqlInd
MJG2rItudmmQqOLtySzj0J/PrwUYkKaCOb22z+QVI+0+TWMQfPeuCPP4iIMFt95S
dQMIagA39gANy9Wti/FKANZYkbUG+znJqFOOsfxhQkWFeYD+VXOooKcfEnpfMlyQ
QhxfgEoG/ZgmIVoRkxKProLKdfJUe6Z1zDeExyf5mW2N1aSDldL3Pn0zkomLxq+4
kVRkGoXUB9NcYLBK3TWam/LyxleHTMyEHZPJ2AJhjxXlqAMjEGceTBzmvQkZ9lxI
M+jBVDPw4RQQ6wd25ex0ZQBz7tfgFN4xJWrt9vAss54slQBHyMtujjcj1xOJKnXt
27b7hkQwxM7q1tdtkTVudy4HCM+GBRKmm+oBfDhkJKW97zkjo4dD38b/KB5ixVbJ
h5j8eimYj8G0ElidWLIHrJT3Pi+e+dUJfKessOtdekL6ETPUztTu6VxXhbQTk0SX
76+OKzyBSVm3NtYQN2DR/BawxrQI5s2rfLu/+OV+o+bmgxDlbSAAjO8aTX/Dyrbb
5snU0xNXIn493dUAeTEZrJ9+Axl9VIf+QwuOYieAbTaU5KlNqvg6Ms7JvIj/+sZr
/QvjwmebxJD+QiK3DWVBhNyD6Gp5ydsPW667jMSPFPkUzQBGGiXe5fxZqZ0I1rgb
jaK+Zl+cPUzalpsHfKdDatg9iyiPf0rIIoOZAvI/A6y3Xoir0gPu/xJ8auYJ0t6K
B5cuDh+htBv+fPo9/xECHyHhJ9FLc0C6z8KaGFdUlJI=
//pragma protect end_data_block
//pragma protect digest_block
/b9epKqb8XKCO94J/FdqJ+ZjFtM=
//pragma protect end_digest_block
//pragma protect end_protected
