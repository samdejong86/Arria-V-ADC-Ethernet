// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H=-!G140%L&?(0N3*6>1_Y@X?)?D,53%08)2>)NBI.WW(MV@V*)B<%@  
H;]E?O),2S6J[E=W*E*P4WNQ*([[UTD[MI\<^CQK0[(@KDKUE'NA(#P  
H7B,W1SS2-5@]!LDXNB@PXH:P3Q:'X6G5/NG!(6OWW!-$0"W7X,E('@  
H)"'!_E7X$RRXG,)B98/SK3(>UST(SV6P,#D27F8#E+SW=]3*O^.@F@  
HF:<M;KLFKF77=%CMGNI16%$_R3Z6]]ZG>+E1LJ53D&/,^F@<A7E^70  
`pragma protect encoding=(enctype="uuencode",bytes=3728        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@R>;VE%QE=KA:-:.H3[(=91062OWX(U)1?^#(^,6TTB  
@=3>K4*O^.962,,-._GN^W'6=H0H+,_56802WYZWS\M  
@B_!8QW\;EI]$FTTNE&S2KH&&BW7I(6;RL,5%[(9?/]P 
@9@XU*FKZZ^*IJ+H/OP"Z@\HXOXTAT$QQ"RUC#;1@59  
@#/$KEXQ]]#_)R(%4W:N_2.E\Q(\?#O8&N2"--^Y=(), 
@)4TR.WTF_OW*"54#IIDO4PC0O>2-4&J3$.IVV[(!>CL 
@WR^LR@'U7BRH38,FVP]82PX90H)$/&N]5Z*]]^!H%UD 
@%@&B-7AXS=2M\.$[K1<;)*;-D2MI6>U>@ QT1<-J9%P 
@DFJ^GI$2K(40K#5.RVZV\+#IR3J=/\7-H2##C^FCVK< 
@B1\".S9XZ->K_D?M>D?77Y.E8]+QW_V'JC0S."$5TF< 
@95@\Z%5<E,_1@3"X$_5C7C,T;1=KXBM]CF#EEZJ#J#( 
@D5Q]2S"(#E\]^=I<T(K]K$=,@G%5,+KWW9VXW#( UP@ 
@P&ZJ 2<C>-DT1A+J2:^=,^5]>KYM%"[!%$&CI[G)R%< 
@AK[1'Z]$ABT5L&ZC"DE*M>YB $ Y=8>Q8ZD-S/98O>@ 
@9IJY2Y&+/A96QI9F\M_9N($,(-[[+Q?1'(Z2K&JW.FD 
@(LB)6V"#D(K#4#]^PH0+*+Y12JY%C"KD">3[M\\AV 8 
@MB7&<P$FX=<E^LXG2:NDIUS0YZGY!2< _1^S>N@&M2, 
@F? )IPB:5FW#ZQ72 2/))NB59/349QMB=@>[!@>W2@D 
@MSB3YP-: !$!L*/EE;W3O&NBS HV?1,\^#=/@ )5R;$ 
@/N9)^LNGBG,>6%K)ISW*3%I+Z59.M%#"*JVJ;G3$!M( 
@JP+0I>I*<O';L+NI]-#R1B0S[]_$IZ\DZ58WE=>*,_\ 
@^B*"HR42CDH3$HU+WJR15)7(EB4:#(.U7ME['=>G<SH 
@/T"0U.J<]RQ./6>]'%KJ?SM(;#E-^>J03X=I^=E^AH$ 
@^:/+O=&U>%&GW<9OLWO3J:QD-+C5P@3SF4X1.PO\((@ 
@@BW-YUIY*..CP!7MPRZ1CK&KPAA960M8=J"W$LE:B7L 
@6]#"%97EBH=0!R846<"=^>-TQ51E<X![Z'J#*:CLM5$ 
@X$7TF4ON8V(M7D")-PN%:A.F_#9_',RTAJ+\P::U6QD 
@+4,Z@X+@#S*W$9F'Y/88U+)#6[JVV%:*JAU<;W,_R\@ 
@?2_*76#*81^K&^@<EQ$QQ>G=-CJ%LM6"F=5@0 9U+(( 
@Q*^MCRS >3455\H14WQ_A;G&8*GY:!AGYF:[E?6]7#4 
@.RT"Z%K2)D9WZT1%I+_CHZ7_,,V]QHZS8>-<^,9P\TT 
@5+FMT:W%C-6'#3[T! 1_75,MYE#HF\-54*J,Z"6B2Y, 
@-?\\YZEV?GZ)N!79FPHH2MQ7Y4?>S@4X7#J_H4JXK24 
@O*X','T))322^SJ#MS=^$5S[;# )[[/RG'JV(1G&2*$ 
@[QI=FBRN@JEEX[(SEKDOL?2$P-];D&]U7!]C_)'^CGL 
@(1VA>ZDX=^U?\ !:/,5.Y":#/&7O(-\$H=YHCX[ITRD 
@JY%@OK;#HT\ VT*  0$LA'%/D2543]H'\3M4ZQC4B3X 
@"5Y)V*51*SG^IAY]GJ[?:'2SE[C2R"8^Q/<6Z5UX1L( 
@C=X:J4@..Z2X02$AKY$>,;)N9Y448IR((^\,I0.CXV  
@&<&$HX:.=8#="< 1H%SY^Z@=,Z,BABDA;IHAJU(F-+@ 
@=!U.J_CMU"^LSR:DEE2\[&$@T7(Y.=H+PE,19@NEN,, 
@*C0?@!2Z=QQ3#MKN>$;.%H:E./M=,T9N6TH.!&>!X3@ 
@#0#[K*%N)9>4!F X8#YP/M]8,2M.!Q\5@ PSLZ>ER(H 
@,0B@K.#!MU]$8R]C'DRL&W1EIV>++YJA+UI#,\N BV< 
@/L*HSWL=[RGLKH.H+@,M-^;^MDBZ(D;"EI86W\;*R!T 
@J5D<+X\B;(W=^_@[;Y2%*U32!5]%ID_;D]7+X(FA3%T 
@H.46]0KC1"*,ZP*H'I=$V*(IL)(2VH,"H]96G:?@PR8 
@(, >5:_*+E)F6_3+>I!EPJ]>,FM"SWQ)V8S2N ?^"J\ 
@PP/?Q=,?J&GV!IYP0(<X#5B8R 2\9JH$M?-V._\R^]4 
@I>KBN&6(JW&WN.UW>K9YD@T!9='\Y"%W J'F3YF *KL 
@.F&+I<L$2\:N;X^['?V?'V4%?;)<!1!_TEM?!84@#0( 
@V\L<G=(L>XD_P'.EJ)ND4YNEV=7&&>\?7>R\^&-6/S  
@0[J_4&9+-6+V'$H_SXHM)]27KF+T-B%LN7C^^:--U)H 
@?Y[F,H-%Y8KA2*@[/O52<!><[@1S?UD+>5P9,*VX6*0 
@ F/#]YR2<8O7H&%<I.$?N?E01JFZ<!=B%P\%)9 )K$T 
@V" ]BTN%1IY1*G-*:/0[#!2_:T&WK,.(XX$XCL^LB"$ 
@A!C80)M;4THN_S08Z1QS$*IHN2-<K*^C$$][*V964MD 
@T7@ABE0UW"]Y2O0XY] -K[Z(@0+W2436.=K_ 1O)HWD 
@Z0;VL9,&>0='HI,WTL A;J-BV;!ZR[*PY0_BWY5M@W$ 
@ZJ*1N,VA%QP"B0LJ>!L8_.O3-2TPHV2238B!^Q0ZU@0 
@X>X?I[("6:8Q#3LC+!MHT1+L$9NT?*/.N$DV/@<4@4( 
@]]QOHJ<%*G#5EXT,")=SE7#Y2<L[.%R)??<V,6G*3T$ 
@R7X#F@><-5+2Y.I9\T?[R@)/U^*+EJ?%I.= ZOF!(F$ 
@M*:P#05[@Q]H6TB8FC#%,VJZ^$MS?<D2%DZ-MC)@/(, 
@>?C6/>-D_QWB&L%V:("R-$/0]Y\,?9K(7N'8;S"=:0@ 
@)SRKVRE^OIU^_F>-&)^/^8C4'J7 3!LWE MC"YD^800 
@O8O5,\H;*?78X^='Q3]YF37?/KEUZ8T&7CX:V-,LB4, 
@+YEFDQ;3X;\?=.LK0',;DH L(YW\H;C$=LP;?.M?G]$ 
@*@1,0K0EXK 4I39E\2Y!"5FPY5K!T!0N09*H]0RR-I8 
@'OASW[N8]O5F44B:S?=)*.M?7VTG_E3HY4WOV(1-J$\ 
@4ZYX:ZV@F[=*7_"-KTP(V8=;[Q)TK1K3G>=J?MM[,80 
@*N1GLC.7+[FJ@'N<4C.AO<4]+]E9VGF94D@;6#?[=L4 
@]G; $C <[IPV7S ._E6RW\H3X[U<FEN/0*2MXIT7_M< 
@!S4TH^:Q2;?X 3]E]>^;80*/O-J7&39O[?E U'-1=(8 
@=**)A-JH]NAX^ZS"-="X9FA$^"R)/4\P\/6"YQG/(T< 
@&J0/%H)("54TW2&;5*W:Z565(78NR981XDXZ%]#M\]\ 
@ !@.,ER!6:X,UT!Q-.4Z &'H_<,31R9O"DD"I93I%.  
@["^H"E538(OVIY.EW<=,=:&'ZU:RDI+S@>,]-MG>3=4 
@^BEZ(ZC5.2-TSK1_^4(>/,W[2;PVO!-0F?MX'6*Y%G< 
@_NPN5Q> 4.;=4UMYE2E+[Q_<BL;QQ@5 8;L).A YX-( 
@ENS!?!BOEY">;%$=$,CIG>R;JAEW2XI*9I]W[*F@T@( 
@D+AFZ8WCU%K)3"AU^?2'Z873[1HUM2)6!_[@8N1C^GX 
@L2N0OO5(,+6OY$ *DA+=46,]<+CM8N16WB$PK8W: UT 
@U^RMKJ2.MFM\9%"+5<<QW)M<4L8DM11?WM'H15=4,P0 
@,\T.EG%.;.713-7+F,?Y)F##WS[!N3":8D);?S@]KO8 
@3M@W+YW5_@!@^XZ!OQ;!?4TI^]NVQSV8O:]K&B6LB<L 
@'RM)(KEJ] =]AMA(7L>]FM?'<Q1=#1.7F,."^W0>=8L 
@>7L)^B/)AI$!-$\_:(@H^@&*U# ,G=D6160B6*&)UT@ 
@<=/?E1]#NGY+(0>YF1R=%LUIY1X28HX[AL>PZ\#C=*0 
@_H<1*&Y:X^6?<9=T'GUW,S!TS_(G6?<#A7R@& ;E^@@ 
@7T!1#ESUT7L'-W&?5_<L\,/NJ]%MVH@GX;9@O'.8ECL 
@7]-ZA%@*9&(JI"&0L!H%LSS]TS$EE<GA!'9#FE8_(5L 
@#^"HT00=UY%Q \!;(LQAY]M/5[C=G^@?.HD&-_PV":@ 
@Y3_(PI[UY\QT 0\DA='RPV=:+<%E^$B*C"[D8]S'LX$ 
@#N:>E^T+*.C=,BO/@P#(!+Y6(07E^M3.+#F.R]D7/80 
@.V'70 ;B0N2"YQB#0GHTP/*+>1RA[D)U-$&,QRR)V*T 
@/AV)EZ]-+XQA*P6^E,M<9709BJX/KNFYT.HH^)<:*8T 
@+5'7$7;7,<#"Y4JX%#8^LNLJ7Y"=D("Y2.@;KY64(>4 
@A4BIN(>Q[Z=M.PM,/RKAUL:E>IE'#>*C8WE]5NI[DF8 
@F>,>OQ)Y,[YN@0!HJ]?6]=#*D?I[%,T]1'!9=\L \W\ 
@<BMO24D2TV9L%AL9[0_IM%0T;4!20*"1E(*7=*ILM8T 
@Q$U*T(TY4X5B/L_^&+TQD+.Q)(?YN,Q.1.N!LXE.D\8 
@3 >:-Y[D7P$&A>H1[<Y5\@;_"N'^V+Q#<AU3!5$;\ 0 
@.^+CT&,7O+]GC9 Y-XE Z[,/*_Z>8[/:]],VV(JV*<T 
@+ZE2,C,(G($VY- K]E Z'N'(BH2$-H1<>OC&[-214PP 
@H-:O9T,>U\@@4ER-\XRV=@$1<2/I%0D0M=U/EK^N33D 
@/8ZX7L#S ;NJ"8DJGNS>)Y7#4U=;?+C<=J7U)TX*'K0 
@)+Q!8>LGE,<_5<-&#R'BAU5;NTB-NOOMM@\]$:IU.,H 
@+S17])=1]R<S:.,!*;,^ 9GG<N[SQA0/!=H?W)TCFAL 
@Z(6:O%D&-#V&S,_F,DO][F8H7(JI)3:R9CXQ27QV.8T 
@^ 6@['><N@RO;T$9?=F*&^XN%6U#F6KJ$MFH4@,<O=X 
@^="WIV&AJ>Q"/P3]D!1$ZVP8;#P+R8D$6^\?.S/"[P  
@13?*%J\LW)T>#*U/7^+FBJE=)(J\D358,7Y6,T>/OC< 
@V0J@T!;LPU)'94VUV.8WK&''T(FENA:8;2GSS++ F]X 
@,00-@(IAMRY+8,S4PC]3QI'I36T9_WR>J1& W<6+6W\ 
@,OTUY&==OF6SSR+97:7<7S:QRHJ$=<X<DR;VYU]LDBP 
0+(%V20[4\V!!K(RZJ4@TV0  
`pragma protect end_protected
