// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Mon Oct 24 23:44:22 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nR6Wy68AHyBpmT6SK0upBUOyqYvLRBLnhOSt2aCXpHZRFax9IsQ7Mdsf2Li+3Zge
/IUAgYRIjXbG49+cK8vXH2rBPU8W/drHDAWm41lH6sx3OqKQeV39d/Qmfev5qpGq
HE91F2fjARnVBV9EQxNA+UQ2IccpBzFCWlHpvOV2+Os=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5184)
vIvlykw3UXqJSf+sGYKxUHy1BgnItGFNINCLM8LEWwEItGQ9Xm1aYQhKfTWkYSU/
iWfsMf3j7gsWaXE7c6auoA7hddqViA5w7EiWzyUwAYwrnsoHYUeCEBukQZroxtFP
brxx6I5uwnqQvSQooXgyRzJkEmBL+MMPvfCZw19rXaE44lu8E13NPbC30muYhIEL
QXIbk7STeOt6hNeOJW4wW4lMQwHWCOGwkL3OCYZ/T/sKQgoZdF6SMZVT294W40zz
1u1JfDfwUFtqgd22moKKoSAGyRNAp+Qmo8Oiz0kfuxvzDV7vnGGGtq14USEPxVZE
OOR5RHVHIddFY9YrJeC0lTzD94iA2nBTf/V7L2WNdy8BGT+45SshmMz8cfr+ZHWS
Ab+pdVQKAla5IsP+OagpQH73lnyUtJp/xq4UOu0PdJteKVdZGC5WNl39JKFYdJyX
nsyKRdI9FhIXoOPeJWvQ3q7xr3QYZ3NP9mPDf5ji1y8BzSzbwkUVUCElI84klIiY
JGsdqvlR0DZC1WRq7/y+4VCB2tYClMSdb+gwMy7a2QnaI5N1oo8coPqPtx9/oeGS
yluhV6AO6oLHTybPXyw6j6fR3nmcJVgEjiNJAi2aawg30fjIMG5AcX1JH7U2hbWa
JSdn9zEuRmxq8uegpehZXhdbkBoXalVeMKB4IjuLQLhkZ36yAGEfH4agtlbmwk/s
FByWJsgwL23wQyIPjR96mNrOIZyGTt8yx8A2Q97b32fHiPLVvOGk7iurHhOPEUyA
hO7qsG7cl1SAyZp6jbQBAT23ZHRUXxExOVP0XNNFdJdsDdyN6ynV0tGzgiBBS/8Y
Hqx95paQjuPbDo5QVjHwMRZJIAZYhVcLTmsgR+o8hdvOYKv1p5hXKWfqZb96yUQw
WDglgXjl4nxl/K2pYrA8Dwe+tjdE2iX5R8VBjvFvJZ6RCoLZB9RBalYoToa2D3Iv
cdHYO0ouoMhydLE87TPrZN7zFVkvUCUOiDtcxUbeYtzOPpDEq7PJIqh75WAfDKmI
PorOZOwQvaBKYFQqNai8CYxAVQ5sNtjS4UE5zck8ObOom0ZKZh+aiYQmdk4g5bdN
xfZ0L+fGelJ1yZ3v8raYduX5cL6s6fH4mLRHQDYdOX2MYcotW2Sg5IMznTcvF3+v
jtYZoj1mq+iy4OHBrXQMOPk3BONoS2CgJ8d/jFwR7IJVNFgnQ4QM36D/yd5kax6U
sqPuKiNqx45fwdKcmMoW15TgXHZ4lUd0DN6Cs1D9EstbDNgPn/B3Wj78iIrh7xMR
6IA8zdeE5WbhHKE/M6OuUqofW3nV3J2SGKY8eKRcFNlHOZLlPCNforwVTZzyJrFq
YqY82py4jV3sRTHPdt93bHLUbBU5Q2Po/AYylOY3pNkP2frBVprm9m/EVHLGKmt1
Ww0kcUf2Lrme4atloacpY8xAnDGztg21s0JuvwMeOiVFrS+dwuCwvZom0vC/UK5Z
dTSHOat+gJGbJaOR4m7vvT4zSst+I3akfkMa/LzEYtmQ+mgoiUL+nbWzlWqr6m1Z
EBybDNgBoJ95lQwxUoZLq/UR3oDoy4cYAV/0DL/L9aTN4D5aB5pG302Y/CpZftRU
whOPwrrn2AytsKGW+85YlXF3WxTbTz1Wg+NfEgIriDPNWVXxFu+JnzM4o4rWqC9l
vQYBhDUzYyc9+dixeZs1mFQBvfwyUhwyUBGykZ5G74kKqNiunoHE9iV8fYQSWZf1
vwwvB2HPH1Au0TYLfrzj8cHxwUOtbXtZk3gQlLhZ5nTEtuK4AckbhaW4OTL3Gnw4
nrYjbmiBJlwxJyHwxKSABgdYwDtVM4/ujdNC5hKg7DOMm1BRkkTPvuAYK8SChvoG
lmAU+sVGggjV5K4KfpCc8nirOQLuwS8pHdNK/tZBkZKN2R05EY0pVhyrMIqvlPSa
MjLvk06S15mw3ZhPG6i9xiY88MxPXqZg32kSfGJ8etSOzT17+1S5RxqMq9onimrv
321UxquouQ82vzsYKlRZ5EM/S5CbOs4oW4eiR0j6edr/m9LDQlCHWht1K3yjEV2B
/mojG2KBH6i3sczOl/oEC3pv4qw+1y/bSNBFbeL3l3HMmd5I36XJ1A0dwJw/u7j3
O1KjYVhbBmtUSCYtqIfkkQHxbObUBYjhl9RmoSJ1N79R2+CY0WvD/WMGqUamTJcO
DpY/HQRjqB0LIXhRQggBq97nSDMuUfybZ8YvYh1WB3J4yuVMZWxqYk0/o3lPu43s
NamwwroTllhNfh24tagYMh6p710YL6KttuGoZ20r86rr4HUAfW2fafGE9X/G2LBk
9m6Io6VrwVWiC9Z1NNAJr4jT56BjfbiM2O3Fj7GdYXyo/N+V9zmkIcRwnFkugsId
d+/7ayqNnmgeScAmHWTLeUbvDY0wcUewkNvogZgNgvj0VNkOTSYECSaJMC7CfJ4S
DY49Q8ko2Cnc4tzxGKeR29TOT9hwD5HywvIPiNIswOhWZvxcJPKk+m4n3YMOux5x
6Kd3k51GUA/+W9zpBZb+5R8YUIQc2Lb2xpX90DPxEqkURy0hSVop2yCeQjOlW/9O
D+HxmZmguE7o91je/wClLx9HJw1g4jkqiJvjYoZjlY50/U64H5h1sKujvPAVfRRE
e6E9s0+pQS9aT8ptEGOgZSlV9qg6oNmh6JQVmUqFkM6bHRAYss5hn+FygRoIhqHE
UUlFT+vLkwWghLtj5aDzJTZyhz96ixnjFqAi9P5WmfoSQoEVo9wd2/kcceGocGW2
LEF5XlLJHor2IB4dbQpG7Low86Va+lo+AQVcrS2zyXkvCV/eikohsl/gbXke3iWo
SLUyKisxhlJ88hQsMcx3rmpzcsNPK24BYuXAyql07OiDyuqaa+WafB+mIBW21YRj
V7viIFxYMupMjBIKqIkRruDv1cTH+Zouzgm7Z3Ok1mkpJMwiRXc2UM6m+Ye0oNJM
MFPO5oZianlDKSlJ9DSK3p8PElLt3kZjdZeLkjib2iB3EVBUelSw2insWITF/yww
Nl6X+/qLprWMUxdfIvQDDgLZxTYBg+VkXgnTWgytLxVApTDUjRQihKVY8KfxW2v2
pttodG5ciD88yyUAHejzzVAZ7s/dvnjVKgA+ZXtv6F/m9uU+WQqPRB1BRdVjepYQ
GZnzS6cBDkh7jL5R3eUO0PzVgDuE+4/q5RRlfhtWHQQFBO0JVnZF4+xFvnoW+2hU
EeF8wfYVAa625WdllcMYk/1TveQCOUNFOh7ySfDOsn1sDlGhz2Go8svWf5pNPNpq
FFkhzizSr6mQ2ZxF159MUngtqvOarcASfqfVcO13KqwrppJEHEU40tSRF1bqXlGE
W9Nmov6e6RE7y5NGdNpFKsE02EifwxsxvICVLZZdSygLpeDODjMNrI0bq8PrZjmf
XhV36owVJOU8JXL+F51r1lhjPkPiCIxZWMaljltaegIEiFTdInXbJzBbzaL9N7//
bhMMWeiVAi1UM2FqLyaIehatuPK52uKdJ3M9mganUf5NH+lO4UgEcPdQPV8QxFx4
fWjmu9DSfz/hANDyr87zhZ3Pj7C/tUxX4z2GJHSBw9w0Sb+wsBNhJywf/elOAYDU
Ruc2bJwMTzgCSa7pbH1FMTjjgq5p/a/3P4ZV+CAJhwZ9TyKrlu9MtjOXBYJhUP7z
pbPLOrLexZx0yCEpeKpgbXrf6YQcy6F8W9aypaRj3c388bjMPKqbcMEEp7xLJHwv
AAGwgf9PSjaJAbsX/zW8Qgrt0mflUr0ohMff1K5GKZpfGfWTQV9pNiKR2nLAIYp6
LcT6Z606EvgMhMO2EiAiTYIRn5HHEcws0jHcLogpidn5VL6ibktqa8fqMTDIr46u
nOMa3YLNO8mF9+82bf6nHrkyU0u0tj1u877rB2rpW0hV2IfAM3z3ZK/zhXH2d2xh
HgAEzJ05j6hRU24rNHUVNs7EDWTP7kxFJyiaCnKpgV64Q+OgeCdd7ieygo/BmL6r
fMsxI8L966r3ZdLPZVfxr0Pgt6SCCRr0xJU/9R+ctckSL4PUSuHscUZMP9MhKSVb
jJ7ciWLGrhCRYN8lqWu8NLD0jWOCM4LX1PgWhO/Ub29Rb9jrG5TpHcA3XaNArvfN
7QYBww4UiPKYZvd/BVLYmR2Mb5A8VC0nySlF/ReCWSmqIne5zI1D0UJqwiR7JQXe
UG6dsAw4RTKONxMv023VQvwVSRxrDT63kc+1KZ/n+N/cUTQ0qGcvn9OoSkT7ZsOz
6dIAAA8u5SEuoi/AMtT5AKSG3T2ezGg46MYcfTuZcGhmohz5M89mjCWxUhXJ39VR
I7lX4WzB1mAEWH0XUhGTB3Fg8QV9AM0gCe8MNnYhdKp1j4M1IgCaD+VuQ+0fKZPA
Zt28xSQtSp98pixNiVCcuQO29nOmLtePalUone7vM5e45OXwQgvtpoXezt/tcci3
dK9LWUOpToMckDihK+ctjdOSZJM0jIygBeNa7p7ZBIH1SW/xpMhvAtc6oHt0qCpH
plxQ2RcgscRriRtNvG95diWRkon8Bfcd2HyOmuoM77W4zl5vr2v9Cg/3inIE3GWi
fj8VIN+f8dMMXa0MfgsZ1jWFyYg4h41nC1JJNkTd3NQMuNqewq0RuwgrbFV57+EY
JM9/3/DD1U8B2SoOImN/ZdpPGWHDq5KhYD5gGPMg/tdGu5Y0r7PYOBh3Hs1YDUae
LmwxGqrn1p/TXdYhRRtDEoaEEydU9UkbNWkR2UnVqdeiAu/0AYnncooelh8f2gcr
naMIVuVRejvLUMNliWindOiKikxl4ktD/hiyVCrkqlJolJAKERNrxIR08XzUCriy
kLFL4TFu3N3MAUymcrv1ZkmnTBT24uNTasgAc5ATrUgAkIWlffR6Ae4cR9oU2iAt
U1YIfl4GF58QcEBoqNrY1ZkieHk1Hub4ZpHRGPjYqNZx6VYqigZztA7EHI5S+SJi
+EkoSMn29FvPFvIykfSK+vRjPjKrrPwz3zAKwh/welrW5mzK8DlJbugR5smG0Hjo
MTJ+jRzHVgkIvLNG9KniucWT7/519u+G51bF0swSubAptdqD4zb1PaAbceUYRIFd
Lg8wKAO2HDmtYtV/TT8dR7rlS0pjTxodUNxlG1+bJvu6znSTXR/yKAVwMP6BoNNk
XvI9iGQVTk4fGVERef6oDbc9siY6RudCcbTUOEu9OeTFUjMw/VnyA+FIo+U05Rfl
fIaczdKzAz4TYySHvqJL0doFol/QrPx0NECrdewPLjUxuAfuAIwqdf/GgFj4RgWp
Tzmd5EMxJHxtFSj3emvifnQ9mdsPO0FzK8RX6u+XLJSphGFX6Quhx4Dn/egHfxE1
ynG767j4BEsLI2Sa9FCr38wfxqYj8AvxQJczAJTmWFAdbKZn1dF84Dur5t7QuXDq
NvGYKvT3d8iR61UO1fwhoVk+2AiYnbRDfpAm7YZSapmcKHFSLrH3yeoQSWXF9Nga
Fg4Uwvn92GKiaROO7ulEbknBaZSzW6Srd8P46gKarTAN8tYd/eLZofX9zsFSWsAi
CT3wOd4wVB4VwvZuGushvNuXV0AHBywIbFtlhiUBKPbsTGeV7TCy3MpP3d8S/IOp
dCuhMIht3LnWHuJUksJSf4oouhuH1bwlRRupFAdJFqL9R+rMEjPeXbwIBYWCdPee
4zjGdv4kNF5wb1fZ0gJ7XCM9j68XNr2l36PUl7Ykglgqb14UF051qHlIotp8bjJz
N4v5GS+fmS+UaqiC0zfMhqVVgkBtzsbeiMS4evvct3fqHLlWdNOXC6JhWrsA158b
EogqgJOCRtBViEBCOaRxB0FDf+JNvFSOQU3ZnOlNidMG9FRTbD7A80d5jjJSmb/8
t8enD+JPBNXWoFRGF/otKEEeKf080hMbWLx4grLERjPL6BTya27i5AkE2VD2z9Rk
Inli9EFRsKbyXc2S1f235MpmWUzF13vksmkRufbZijdG3qgkXFKMORP9U7+2xlXr
cH3vbenMMTQm/jPSU7mMX6YHpA2HlVfDFajRQSQ/RF645tiGNEhgCzhUBBlD8zJ0
aRpS5yWoPdt25R9SVuzVN0Jn34KMi8emrT6+B0DbjvsmOXR1+0ak/26QWztX/GAk
9mLZiPJwpXZwDxbmNbFItLm1xnkicJU8uR99BpH9uhBjvanKsRYszHc6b3UYv2/9
6H5Xuwyvlwop2RezYXz2IfAje6NMt2VHspEYXyzt3C4Ugm/WQTvASJF4h11XRfks
JM1JknPWkKIHro3XyaEmYCBwz+nHs82oI7duvoSAc39R96UPRGDG0koUZRpUpplX
CamFgz1UlzkL/JnfEZbKTymybG09C8Y95cB1T97Vw+i2RRAIOZTGC3Qea6hAiS7r
0Gjq5ElOeaXNi+Q/jxVFi4e6ryTu9VB9bbzNd0uHj/YtQI03BOXZ6xrVyA52jg5Y
ztxPDyRuIWTCJAooeB4+Wqfsw4Te0/rVXj8b+7ufegF5uzbp+M+WczEU/X+dpTZu
IfjzgVYpgfblNzi43Jsm2z1bDABfgkAV0XNry7AB9b5PKfoC1ZaUQhWv2OmYhtfc
+20wBZ7+tBsmyoItO856vGJdlSRsad3GIMIl5wqxD9Prwg/016iu4zpK8Bkk2beA
zWePQ6izrBXRb2R59+PzP62RUuTUVR3WOPYR1g43xfmcGZSmAfbPViNE9zNgvHHx
R9YrWpKpBacdEu0OvrSkCDzLZ0Il9Zg8V39s+CqLaFbG5siDXtg2c6cj6v5Nb0hJ
Thzq+mPY7QFAnUr3askzJlpnsoBWjgEs5bN2cC01oQEQX682E29Ij6s1wQ654eT8
S1J/Vekl+fhbTfswNKR92SdqKuGzeapXqkkMu4gcf0pIuzVOxGRbBzzryY6r8W/H
8KMWxfUAu6/+2uZLvcWv+v1NdMDHaS+V+Ct6beAq4rG4XZIsZtqhgfL7qge28ibe
`pragma protect end_protected
