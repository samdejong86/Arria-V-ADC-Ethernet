// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Mon Oct 24 23:44:22 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TCuVMUoVUGRFqFdjlgG2Se9/W+HT37REJhC8jvw9akNcQQJ/qnBpW9p5YEQ8tl0N
0HS1KniHUehSjELvhsX/FSFl4glUFFpDvHOVBZlk6LdWlwDhbA1WjPQUXenrs3VC
y1Er+PinALVasBkMfdaztEZmD+dspJQ38MYInAX1MB4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5696)
2WKVYCqm2/wLrDphWsyPk+SzmAyZbVLhWO2vYMKgncsjwzhlrbu0hjPkugj7Su2J
KgA8QxR//hyITbAnvqp87BxH+SfTFFe+dfx6RS7xO/ml4ebRQ7imXAsuK9Gvc/yM
HbGBh+XVMCNdNFKk+bJnwYaK/dMyV0Yaz/TLmi7gHsUbk2Szfs++t4aYNaN78Lvi
fdOGgGWFQfOjRtxhvUYQXx5xvPVOw0vGJriTn650j5G+ruRQpwLxTOzJn2hGHo/n
81RoE5FCZVbJP0FtTZobmpYpPL6Nlnu9kOKK8ckJks76yrnN/P3oyUEZtHdqvwhR
3CTpaVRw9AMF/ikiQ64PGge3qCN1MgevuQ4rKfSWzhMCyOiKoX4fYafkwCBPAkNi
NHAVMd6J/hkmBKjv8laVJs2rYHO/HJ2v/huPP0kziELlmy9snRS6tGs+cJ6I3J5E
4P16pUREzw2A9lwc0nso6yzmKgh2Dt0F9oA0MMPCRCc2v3QsxQgJEzNoPIWXzPzS
xIwElTHds48CvjRlq70an5XK91x/HT18wnyddXGyTEQiYQbBWBj/bMpiGaTgUfio
V9IzJ7cFrFcSOeBVDF8uQYSL2xtGMwG0bG6TiN4DsDXotTuII/4F2W2l8QFpVOKZ
FZ5ywnDO80Pkx/FioyRS7F0p7N8QYDrVrsoHhyzMaKfgYb9Mb98JSqsFewm0uIKV
LaDJD03vovdEsSpDWhBM6DeYNeGIdcwOHAzbbqfGb3lWUdTcBr/lWyVjMsUqHDo2
cNsKGVhX3Z+pYRVnUwQ3MkUWJHB+YAOH4OMh9XRzHF3w4WarjUWZ/VUYCERQDpnP
xAEOEWuxLngHbuv/qZaMCS/7IXMO6uX9R3eI80BksdhaSJix3O+sGrt+OLGDMKCz
H8RFxHMaBMH1omp5PuXAgmdXcCVE1RpxevkJp52vo3jl7TtYyKn5vga7EIxvBrRR
W5/epRSgPhZffG2S250sa2qZUNevlQamzQkUpgwTYoITPGWWZk68NesLwdbby6of
vc6+9ugM36+D8dguRTWBkXFlptRKxIYul9ieXqJxDHPcrV9jRsHvzavzWJdfB/si
Zg4P7pZEI/7yai3hDzhAXTEduPlKFu3KlLqddpI19Z0eBRynDswrjpkY7UlkqmQA
Jol0nCTfAMkC+fkoHGTZSlphDhdpzQ9dOZEoSx9thyuH0DYxCUz0PvN7fNmFsWYa
A0t8ju9I+2V8IsKkvWkVMNOjnidNtQGEtslbf2ccYaOp7WfI1NFmcwwxdjpl5dLo
x/gAVdTx4j6+gCGdURK23fH5llafR683PIGtLhXqBxksCfSt5dBjxkUIgi4WexEJ
SUUgSUIwlKNGOx8znjLsh/rQJljQemlQfzqH4G5eXhkZr2xUQUB1UZu4WFz4PiE7
yPDEaVqp46AxayRxXbVWlcdJE5py98emY9fqVhqqi5KmmGHi3WHZg9S8hcvmX2Ka
bdpWZkjL7yrezC1/Z0MgegTXL1DYUmS/mwPb5Y1uDaswekXOXbrwaA8FMjGOE+2Z
mdfP3rxbTbjpf2qAQ9VpsHtRAEYs0xir/EiVFSUvSgINtwWrauhCVB5tvlDJvFlS
AloTuyj5RBsaX87+EKsiEIvlz0b2u6RhILnArNVLEPPFaM44i1/NtFm/vLwL4jQB
3FLesPrKsl08aUkxu/Fv6+ZKeqP2we8wZEAI7k/9Shrcit7E/Bioy0T9CXwp+eV0
D5BoqUjTpCDVcWOGHiCQ7wBJufsb9e4FLxKj5o+fxr5wALkkFdbBPGI1Eaws2OWm
NPqwlzscQPjTWtcK2jHR6aaMYFwu9Bt6IRH3I5MbGWgMYYEbPJVdKXdQC/XECYyX
SNY0V987eeEdF6dw/VLD9KAnnSZLii48q77vMXp58JXG/58so1eY2gOy4ZeztAD+
TM/f2XrM+8NpMB8Cp2sQJxUV9DJz6EtScKdEHM08mbGLn95Ly7ZUEvRESbvHHa72
8zfZd870hxfGXFaGbW+snHZ/qyeoQXGBTM/2auJ0kLWKMROOszBCsIsg5GFvvHdG
M9uTvif2khcIIrMPQ2Q/KRxyE6HBIBrd7UX4JDjLtylUTnFD9FNHkZj2Mib9KFsF
mXMH7EgqbBe3wU+XFi5dnj6P3yR3O3cYwGlTf6tVjieDFPAdpfrlI+5XV4GQX2fX
dFvJqqlX8Qqd/RfYv2QmnGWxxoOoGGS8mYfmWsB743vZPgO9I8Db9LPDFhm17Fy4
9Ph4P6kKx7nD23mwPH159hGKQEgX9PQUYA3GvvMfBqsA/1+SLHHEp+1SMJ0sGG0N
/Ig9AugRlD06qpEEei0fhwAYiHDUp2hWUfeFE6znKZjBM5/Blg0eo5vd3bKrYrer
nO5PsJj2wbW7uLWAX65WHv0N4fYJZlLrRp2Uh2W0f6RlSUoE+utxUbxVJPk1JYzx
zkD1tMwGfrv2LSiyPp2oBeyNc7HlDJUQj0CsHHe/3v4HoIpsk6rupEKoKOXQFBxq
NCxvMCYdHhaFDiq0vtNXoVRKav4a/cgvKStz07QXPO6cadocvCN9ljYuIHaBUlqJ
lJ5ctCILApZBuil/ctB3cTmtxkXwECDBJcwomAPTZyrw06C00Uc++SBbECZHARyx
NIoHy4RltWoLo72a0R0QyodWriZcvw161gdxacInH9XPRQEyZgvx6bnc1xYjhPgT
GXShdoLqm2fxNvJgY40SARZK5QJ18/l8SN4w/2AOtwb0VPkoMtk1Z3VHyXtdRPbV
EPl0pNsTyxz5OgtXyrtNiCzW2xxDi/t9HkAWoo0gVKjvo0D31gF4FyeT+3KpadRM
QCuXCy1Uo+oz/WDV1craYsx4qkWFDLM3wjk5tlnbhbOLSgAOxmoD2JvhJdAp2t0q
d1wb/E2L9gkolR/di2Wgvscz5rox8LXmM6AogIFS1RS9lNz8gCzv6nnZOnc1RRtD
Uh16ody0GTyLWHnkj7ChmJ0uJB+6qyO5KrLwTn0U4/Lg1QETrmojEK5D1bJ7ejYN
OX7JkfK+KSID7pGzptUPTR8AL53oPS/OC1inzNfnTVqcMYTo0pttSpipw20U6CT2
ayRLVVeZ2Sd+CdI2upYdWpg3SZEEnAH3BW0257AfaWgCYTFM7J4LDEvn8uVcvcvm
hlSd2ex8OWkpoAPhHptRcKBEgyieWO6tvc1EMO2r2MxDLlDOAGRZ9fWKIdUjQStc
uRp0s5pHfzBmHjmnFcC8Z2YxDkDaa++CW5vgT0qtWf4bDp/Ggzzrhu0VMNQ3iRpf
1w5ZkMxcZChbkDlLicfh3pfZsrPbbapowf+bWprGroVeeGcnpcBcVdR+DAcbHqG4
CcqjVYjCpfd+2mjzbMOnBfhqejhnY7iA7Jg+dZjkDlikruUnS2QqkfDFl7FcLKlA
Z4/fSE87meRM+4F/q6Ot5jkejv2hSEB3xbSYdlEuK22HeZ1unijK/g/fIOIBDOQa
bV0gJXm+kGEZi/6kZXPCqICklrGY3lEG3mNNC10FaNCls9ad4jl2qqDeLX35Zxbx
ZYCTROz3fBzZrh8jTJ1L81fZlmyIfhkAYCzKQEjYvADN/M4UPtLJLVFXE49pSQGI
Cn9PohIt/GC23Ee4JIVpFxcMsjqR4/gDDgNCmHd5Ppa9ooKV8s7EkiiJUTK5mKk9
WqWUzhArAYEb9gTG1KJ5h3la27dtJT2Pbt6yJ1nnLUZMopILoNLFDNwM0AzYPHQe
5Dc9ZcdnVW6DM/l438Mvc1eGYqNqlUfge3uOp1frSUCbx304LGxd4Z6SmkjLsRZ2
nssa5h+D8MRz3HVgJbfkaF2Ae33eJ1B/bhBWCW2DWA6i05cdptWrGn/O6QrjxxdR
eWSPDdLkTpz08hvEloBUzN2XgvXNsPsc2JdkbTm7nwDV34IecuK6pG6/o2w92Sgk
P1lWMzJf7UsEgKz/broWOfl47FDUekm68G2erd4dI6Vi2Q65ugeqrG+ewzqVl9BT
LAbuFgQcGBc2Zr1CP7DK7EuPBPoVlDywE9dOCXE1NQpZ5fN12CagCzRoJh8RXlUY
GHUZDu+toOmIr60y9pOIVCmr7WTjt3G474H+6irsK5RlUh/CTa6TskfH7PiaZFeL
L/X7g1eXiFhFsS4uTnGSvQBr1qIGy6ILKxUeFRFUI/Fk3ZYZb61lnTbUCEGBk480
RpNL/pJgTNIjSSqt9dlW4xdOQGalnVl1zQ66FTO5DsEbDH1sdn0B9A0RXnINTkp0
iuJCGrCiwi9aPGs5jvODf1gb9ECJ4U1otpUQ8O5/A+r3dkRF2tbRgLDpPMXEy0Uk
yoOryZF9kh7ctziZ0YGPvX5fg9xwIav9I3phTQrbWTN0LIAb7X5s9qpG285Sgr3F
haDpVsGudLT4GSsb4n6DF2RiKu5h1OwdN8M4O9PEP0CYOgl3eZ7HOMldfwNHPpIu
W2E9eB8wvStN4ENVrGv3AJ9mqMP5j0b5KvKJ8juyxC8mAnB7pjQM/hIQdlfjLzPd
pMDOLE8P0UKpDrB5o4DmgsHyyq9lfjLQTGmebpKbePDgVhivv7B/BVwUGawW5KVB
XdPfgxo1G9pz3t4WKAF8J0A7Cc+PeN3Ngs0UScOZOASUk0tLGELGEuFD3zD3uxiw
hb42AV5Zd/xyP6PoPXaNLWIRv8o2HpusZ1FkR44FPeSWs/UNHEGoRVN9uH5qfLCy
e16lNZNfaRoGpuhwKvT9mthhvZE3KYHCpcgcBwttI/cn21lu92TiEvsDy3BlmsKW
YJh42V1ovj5CTpVxp9AYTtOrLMFsGr9wW+bCbYk8tXoSjSe/vyoSKZwwgr0Prm5a
foydakU5qGiVYIN/b/v9UkGCUEWHRytF36rffL66Ze6bCcIXupHXySaH0470v/cm
phaLOL/iCKgaJYy4wOpQeJX+uXubYWeACOAZWULBnTKWNtu4Ljxuwa20mWsk3XDS
7hxnGbDG/8o1HQFHkH4Oi1EBK/NYbfnwXTUn3pzjMMkbRFrH5Z2v1ufrE046E6hn
ZOdkUWxFAboKYKBB5YJ8gadEjBu1VFUtjP/mN6vPiGk75eQzsxjnlRe+SPOX1R+h
ZrMwcYkMPVc/1iVxNKLE81DcFeCKfQ5j2Ex8gsSaNFpv+0GU8HO9mIbSGIKAHPXv
5CkDAUBZX3LQizQUsz6DVjLKhMCXaO8cjsvc9hBiqVMiCuuGYdRuvDXLOvyt/4E2
y0GsCvhnxl2btw6MXFOmDERtXdTwgWFALC61W3ePR9WGmQ+fcXsHz0UGV4iCXcJ/
8zFf/gvLDWofw6qYWQ2Dbtyvepr49S6LNRbnXYYFq8c9suVmarycYZ9NoZ3I1MDb
V0HqUWm/Dy4okteFPOfdTwoYxnQ2mue3t8JsGFX+0XeR00f1YCKLsryPrXzVTOxV
MWRskckOEuz1BrMfjvwgkPaQhG8lN82DRonHCqqbUY647ns0ZVzIqsEdziyN5HaK
g3zNPNvPbdL1+MUPgjCw3CZnvLk/JJiKVcX5khnHKXGKhkwBZeNesdC6i3hD0/DE
1tm9gpEgYqnKUva7GyioeYN8DER6dcrHlyfREcWoUC8Zg7eM8+0+M6pG2L9kdpPu
PCZkKD8q2Pm0HN33eNqVLz7KDuMOK/CCIougMd4K0Eq+BwUqGBwFnxQz/CJwG7wb
vEz/TkJ5YiMmxEe+vzN3ZivY4BSylxhhUGT5+ORsqZjUB6VXh/fjfSggT+12O2gb
I6NH4xepzcbqpvGg5FTU9+T1rO1KjAnkbNRx7FA9usdpIDPwMTD+wymCg060eSZc
B33nRV8zafLLIHApOTahT0DeXdxWTB4kYMM7MgRBPvLBhgdNagtEC/5Ppg99bvJM
71JRuvjULiws6z6Rr2x4Sst/qD49wBHUp/P0DHqUUwFJdC7ASCFFH19DbewDbUX/
yWzOucIyNrGUhtjOwJrw5tLu7L3hyGguD+Z8Wet+vYATG1cvZLtN6CI+FJljf19T
c6iJdEc+0oJ5U5CGLAV9yyshoTe/Bnjd47nLxN3MQYLMheNj7YfLjeBBBUba8ZDu
yrUfaXMRUX8EVe+30jhQFzmgKq1jXHr2naITcCzcqSMJ3jae+0S8pLqveogBNeJM
qvq7eJPxN41QNszhsokWql1Qio3MnTdqAcLFCkaC+N3uZ8Dm1ymFa76T0BDp3w8H
Ps1LSgZRg6dQ1Av3asPjI9zu8P0wRNokQSrj/4XnLS84yL96HyD3OCCfXdQTzRgW
HXi+SjzIbyBVot6CrfxOdJ+ax7IC5A8VTQ5gOX57pjmpa1LH1ziIQ4e6M/iU7EkW
qACOtrxGuCFOQLvmsK3L//JAjxeLOt4/KncXxxSoe099NiISMIv43UV/oHSd0p0m
i8sbuHdU408BWBqYvQHwxdVvPUZ9fhWLcaaf7jWXHpClxDLPCbCvSa4keAjNgnGo
wvv6NqpisRnd7NejRPkY042lxNbkvAjXkxWhVRnNQNkzkAKTF+geezQFLCUToLsa
ubUFj33fnqQBNyBZLTrNxcTnKOMQB+hYmrUwuosGmtk68Hbby0pgpCrc5o6d5BwU
Vk9hwSrEdhQiWHTHBwSfttbtMuZPSH1Mv0pUMaShptpaSSS64SE5pMh8kY18xTbW
o5H1bh2Di60kR66OiqTfOb/Pn2ynGDGO9grWxDNvAhQTZnaVX8FDsBsVz6/QvcuO
uOzz/4I5YUpKxtlT4nJCB6X4hBkzL1CJIBPUYh/hmldWusteYrB0pbuj9aIJ3Asu
VP3ZNegnkM0ExkxXoD8/Jhn09SY+8dxTT8tNPGyhBUl5J/42He+2bqLaED6uO9mz
Bo2JMDf/R+OZKhNlBE5JDLhALcs6OQktVxPA6ZGKFAkM2xxlchxpImXnyY2yiJ4M
P6xqXYkE16ZAojmgEAWa7eyY/bazJNd0Qf7LGrLh1nlK+o84Laoe4PZungVPafEa
RdVFtJizCt3ueVS0cU+iYj/oSyHYtuzo065Tk7zOWlGaglGj4KA56sVgwFvKgo7E
2p9pKIRMF7oLMv2kC/3KgwXiKaF3zGncEF7NUOMewZfhLQqrN9nDURD8dBbGtEC+
AFP7/d5DRWCrs+Bgm2Bl89dP8hLPbJuy1nOTpoW7IIhvTzZVTp08nTTqHYjXl6N1
AYJtJbG2ZOZzTEbDzF31J2Q3TRdMBZYwIFPhwzzXoH4BQTBV14ZQtcx1XRXcShAA
lYShy0G0a66VG83xdse/Z5uJ8bTFrnL4CgPCZUerJG28BbShNiZVTFOnX3KVamjr
e3oDwgePAAYQH9nnLqykGrx0FvZEx3Ukl9c3/uEyTWNwRBUCx3oxWGgdpkg4aAeW
A308NCpnWALi+zis+bekw30+OTJEpF35gS+b+riTfadeiOSZLZ5h9nEqug/Y++rt
WRohnUBYg6Zy/1EMHBHjeJhycEHUY0R05QzxU31fDH4qd0EBVNgZFRQNNKRF+qw8
tdSRlGLQuclaXqSuU8DVc1Pg4IRvEN+6H/QrOuHkum4mdzJWaWzcApsxXlbTiFzx
HEcd380vlLGBBHNlatnlaurTfheH6wU0PC1WYzuFyCaNPc/ATt41rk1XbT/wUIpL
+vH0xreVgEF7U5nLkyHf2P4LSwvuMPkhI8IIzDMoqLk=
`pragma protect end_protected
