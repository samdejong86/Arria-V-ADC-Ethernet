// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HA9%!;^B*V_46WE@3IJ%',=/(0/$3.1G3G=(:JX#X*?>[_9!N8[KB6   
H*7741[J8[=8@0NT"5DTN?IQQ@*L%P9OQL:WH#E'HY1^K%O, *HJ.ZP  
H%=H2:>!(&*N,*R@.D1\([VR-_BGO7"A),>>3)CH@Z,PFNR0[=9]0 @  
H?EDN@SB%'<]"BD8 ^F)+'RZA3R4+W=OMHNF>"LR=$#VC[<K6$;/(X@  
HTM0\>D1*<KX.6;Z-E%-7Q_3[CZUI6H<@S7+ZDS<JD&=5_R-C+! ..0  
`pragma protect encoding=(enctype="uuencode",bytes=4464        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@-A9S]GQJMG\D8R<U9=R''>>P[D##TYO0OP89[?DPJZ@ 
@>EPIA]JJHQ104W-'EQ1?89 ZVR+R1<8V %\!5L'1C#, 
@!\G+?G;3@])6I(F,9LJB_T67S6_.J!6O@;H0YWHU72T 
@KK \C]=<)]T'X;W5093'<@5YZW_%K*4R%22L#M^BL:X 
@1218.R+!:XNCW%%5N0>L[>)K!EF,P-<V$KN)II_S\1H 
@8Z!56Y90'#X2R X-8#ZR2.%)%8AQ,2R@$7\Z0P]^N:, 
@: :G_]^O<9I%C>^@3TW>%N3%%4';D]CD%U939HPUFN, 
@#UQB/5=9SG*KU/2*J>I_F5]PM0RI]X\Y.M= (VG/TML 
@@CM.1NS8LLG:Z3)K"'62Q>NWIN>NO&-G_D38P[>@1)< 
@+J3:^?BJBP\ZD?+O2RRB&UO;!@6 $& &[ZOUSUORLR\ 
@<@%YK@K">@UGW[!!41AS=H5*X[X*I[O5)XX*K[ \U#  
@,^#"0-)2:-T65+8MA[ZEV8RIC0/8S)OG5XLGGFQXJTD 
@Z<+3^;KT(T.''3%H3]D&UVQ63:TS+/Q"+PW%*U5-0O4 
@)&K,E74C?$_20P82992.)ZXLJ!9':>!2AO.GRSYF=D\ 
@6@>57M-[2Z?XR'R)/FDTR1@V]WD=Y&^B6O\^:[;R/7H 
@:QX]+:(\^0@>CHP6$B!).+6[WNC=-@+7R89M \8MS>$ 
@-*TS6_-J[BK95K:A5ELX@(4/?HXI7>+%7NH#@>=0!), 
@<^&^ET49/#"?= LA(L@Y);+ ^O;/MKC:)T,-8A/^8LH 
@X)N_%%'>- N!/^!WLR?5"@TE L4S"!C!7WFX3"10L;P 
@LFE6F,6!17[[@+6&R$IJ:25B5WM<]@8ET$P A!SQJ\L 
@M[(HC$GS5Q!(JW .!"7(1SQX@[KST!LL.8]5YB7TM,0 
@JK*+>_OM[?HBA/'T6IBU\ +<"'=K2(L[60,Q!K_&YV( 
@G(/^V1<+WD,D/3/,:U!"=<>D64UFGD?UJ(V8B[9[)4H 
@1=42^VO;#K"-@F@)VAEUSCMS6*9K[G%GV?<ZK\4*4OH 
@&C%@PGQV22(\D0[G0#R!^!V6X%:O701,]>\&#YU/MZ8 
@+L>QL8?^_I0+2J$"3>TZ^?I=R_*X4%EJ$'=2:/VR3$< 
@<W#-HC>Y0?;=:YT4G($S^C/E*90O#1H[P611V_MRH=D 
@>UB(52E%9,1/$\JNQ<J1ABZNC$MP]I*5Z6(7:)KN(*T 
@SYZZ'W@+;D-GZ\L)Q!W$0Q4S"?)T=^_@^K!O>9X;&<D 
@7O2%&>_<KDG3=+>I+3?WH \-3X16]@6-GS&C02JU\>( 
@WD$?H(9%7"EH8.5R=%K-B_25EU2\)&<F9$-?!"O[^GP 
@?1XF #0W0KK;73JC'?&\^VB(&4P#CR"AC9A2."/3X>, 
@I@)M]J-MNQ,),AK&HTN#J?R?]#]J #*@!)G/C\_=[/4 
@#7JZB@!6>IR#)PR062;\(<5YA/HA0;N@VP+J\#:R>*@ 
@7+G'C,\) NAM<-S^,O3SO44:"_C$:I[CU@C>,'$O+#D 
@HULNT[9IM.$(*LB;BEPV$Y"D\S]*1TV'ZQ/9LQWD#6L 
@?N+VV$IM>WP+1Q!0?0"-%7Z'$M>K"(&@RI+<_\XUW/0 
@A7A'.]WU0!F&WY%V=/O*U7!PZJ@Y/E>!ZV$$-O5]IQ$ 
@YR05JM; -HC@CO'ZB5>QS=ANP07L/Q1)2?6D]5/3&]H 
@;%+9CEGZK'_V#!*%6G$7>29C:;31Z)*%WG)[0;@30Z( 
@ '79F4ZVM*"A4*IGT[O0FB8HZ2H3Q14/B-YFL/2ZDR8 
@S*NDC@):Z'"<0=#!QA#TP['0(B9<8-J8VK4V;N70048 
@]*%'6J/]A")F(NC'D?:.2*/Q#E9H4'H6[)WKHP>[CT\ 
@']2S&%"Y(<?%QA2PQ?9Y 2'=@YSXI$NC$J,E5@CLFT< 
@J Z9NNCP:$PPK"G9I=-G%N"A#6S,QU",.]!BHJ-/6.0 
@)0GYGJ!B>_B>'?NKAL41TR1[^]Z/RBH=;W@+=L(RG74 
@)SE/SB!Q8)AY/3P!V6I00KL\XXRT.+0<]J+!+K.I\O@ 
@XQH3S9%F0B 3NV?,>ST?O @>"&WG]: 32$'1H%:YYGT 
@27W0VO[9EW**;!6Z7]6ESF*.^VLRG[/QO\TJ8.LK[38 
@>V.\7^A@H4\7EOX@_R34ECH4+E(Y'YJ4&>3-KF^D_P( 
@SK4/*3QU9N(UM*\Y@QM+B7?#5JOV4NV.PD#Y /6[/.( 
@?5Z:PD_@AIJ/CN-2RY$0(CGR-9MC@2;J)!VH\^[GPVD 
@&9O2B:Z0IO]VLTHJD6M_P\*\US0C@Y5+X:';2(?) T< 
@FY39EO^A$+G?F(!8S4_WN8!+=#EH7W4A5M]&31JF<L  
@]S\"/1"41>9S3_FEM^NAU&Q^1#I'.6"FLK8XV3A/';  
@(H%?&A_XYK6+H6G[J<Q)X2=D@=45"THR[%R9(0-?!_$ 
@D/:NZGND'51#FX),95W2Z K=NH?3H RK0^C._( @4SD 
@64-0XS._"0$<SD9%XJF"'_?5]AA:O<9&$^Z'MTZI&D( 
@*O9[P$QL/WB;;XRUTBFCS.,45?,W\_^B\,A]%: ]/DH 
@]TR!WI1! !'@K%&Y^$$;[WFXE4?T]<84CM9I'"/6Y'< 
@O$+*@@=BL$!S>T/;*;N<&E'V6. V_6AIH?K)IH'IAL( 
@8H(79]8O6#C3D!JB?_WC"3D!S?#M=:^=>X#6G*F :Q4 
@2[B0YXN_"%*()B[ O5G5%"G7EC/?UA,.6XNR&(*-O.$ 
@VZ+0 >0BD8,X#+$$?9#" I;!D>%;T^T(W[M]C?909C@ 
@ZL5(J85W4?W1L!->N=[]-J7P(CCSVWA<":*J/FGTX<@ 
@]A9IZNNDW&:=IRHV?2=7%.JTU*3!P7X2L;>-^SU=Q*  
@I]TH9,X$ZTEU1GA9/(!.I6%_*RZ,P!'#\>GH8FU#*R@ 
@61]M^S;ZH9X&.=&Y^=!Z)^_\ETPA78)A:'M]OSP3.V, 
@W\;J*/-P309;MV&A6V&]D71SRJ]&\,9^)X(:O3?C\]T 
@]9"N;S$"/CT\)<]H=+20@/F00\9%S#T&& P[NDH2:!P 
@L<<!U+<>%"Z)+JDDAS_+6'.*5A^\^W3V  Z;%Q]>L3  
@3TRE__\A[3*T4Q_4C3\ZF0Y::0]4\!Q!' 6<J]R#J?0 
@D5*GP09AYX0^R> YKS;&<N1:AYP)OF_"C/?^%ZC7* H 
@W0BD.RE'H!7PP](:/AS%6/2"6"#>"T2C"M\OLD93=^$ 
@]L]-[H\$/-1##8Q957 *J+6[N>L6^7J^=!-W?X#X0;  
@Q.B#29@*V-:'>HY15F>PDW(67RT@&1O<8,([.%*0NR( 
@S!^LY!\K^D+"8[D;;S_6YWUP% %;WE2C+GK[WM8QKEX 
@_QW-4[2V96L8KXFMYQG/$[>_IH@5*?-B=^TV4!<VAV< 
@K?)A>N*LQ/JHV$#D_.)WC^(^=#?8-6P%ISZDR@)A:Q< 
@")"--#HT XL]'I7 GS\COT7TZ%_C(E94B*;.RU_*+7\ 
@MKZF>#YVY"KSS4H/<7"<NF:*#SQ%KH328GL[-A*.NKX 
@\]D@]!8D!.8W>*W:U31I6\LAK%VJ$U"7^C_Y$RX_+.P 
@GYYDTJH(_?B_ 3-.&>TU?.>DXO[^^T'A0XS@NN4^%F< 
@?3RQ>0F$<K$4)#9-$\^03<F(=#T??]41OI;7O*;9^2D 
@=39"[9?3$">#8#CH]6E/! E@WD>D9V R3=OCFPBMPZ0 
@B40 [4]U93*%_>RH5%!Z_VU-U!0PPCQEWU*'602S$Q\ 
@J/@<ZJ7E\\0336R'2,;I@8!V3 */(*S$V!!Y0"H!IQH 
@+F$EYFWYK-?=2DD9]3>(8NP"L)3W+1W'%ZS!%G!R+'L 
@OTBSJDF-S)8?Z&Q^4./%)A2_K1#&W/RT;"5!$8(I2'P 
@T41<*Z#:?B04.X='Z,U L4.D=0UQJU8T9@RCN%S-$S( 
@2S"8 I%_UR($60:+)T;Z7%0N9[H/,M>T']_3VB"5(8< 
@-ZG,RH(8N01-.2*1*F &:$A^0_^GI9/&GW)EP3SIJV< 
@)_FA?9AZ3_UBC.N$OQ2E>N34D_>KM'_JU'Y\34GX4\4 
@Q"5W#U&L.)S.5@W8K!]N)J>U;NELS+):'D2W"M1Q>-< 
@(J;20&9(XQ X0SVL@;,^/SK4Q:=4L76&FZG'T?\4(SP 
@^Z-ER*IU<Z2\X7D7H%"'(J&%Z+E,@576I1."O2;,"L( 
@9[\4]][$7LMV<28Y"LITY+W=/E:.5KZ04^@6TTP+\7, 
@]/E/;*"4L"]Z?D*]9(X@M89N2Y@^ONIV4CR1#),DU)$ 
@YZ+K=NL-.U;R8*CQHL.Z7LY@5!CVAW? HI='IM,,Z[4 
@^ME0/V.N@=[U7/A]CL&N*_UXZ19Q?1O 6V.-U<IGE:0 
@I&2S3#B?F*2?A0&(![ [ <3AU.S=.I^QGKF-1 ;JU0X 
@NSM*+D3J*PY01/41"(J_1A@^?OXJZK<*#KH7$7/]XP\ 
@^K5)>XE-$XYTA_4QS\/R75[TF8").NZL'<-=I%"(1PD 
@\#8MJ95O, @N?AEQ@ J)PYWP<D]+%== 2:]C&K"HF+X 
@-EVP;; >'LD)YAI#XLLEAZ1HTD4VUFT=8F&E^F+A&F@ 
@2&!"CE\OO+>]J98BZ!9@L/1EG;X=74+4%]8^EW>2X]\ 
@$C=X4Z_#V@MO_@$ LUH>"/5UF+T.QL%D"JO'4'X;$\4 
@Y9^G8JYI1R2KI^V*H%3/Q05<[*QS\ZMN>^#FC:['Q@4 
@VLT"MV]M+J@,#[!_&*R,KC;HK-*J?=_%@DBI@!3 :9H 
@*EBV4R:.0V/0KQ" Z'#%!@1AU@R49.J7-T^\"C9KSC$ 
@[AVH<;X+?*%-H6TE!S*0'=C[Y \:0&P+#'K =9==45T 
@]/Z]*?M,*B33"N8Q1:]EM?T(!@I,NB2"6F7M0Q 8-MX 
@[W^&)S3<334ZT;>L'E#4,RB^MV)B4E(F11&>?6>43J\ 
@(7Z,9!K1-82H[YQ\)<7LCQN3[6O0LB*OLI; 8OWO"A4 
@SE-K8'[U8;"X)*?#@O@HG<K%_(:^D*8,T2UJ+(,958< 
@CSR >WZ<? ,-AB$$P+2H_FF+8)(8+TRTI7OB<;K)8NH 
@NS,U(UOI@I>_+#@(-'+G56WG+>LYC;/A*P/VG43.U+X 
@JW,O>-1[=2BW3A]F=V<P=MVNT/<QP@Z08ZBK!$Z?-O4 
@E:C]6EG1JA<J<],\B>=@2#_ N%K!9_0(C$ U8)WC,<P 
@P3.-3]3>'RT[4N:*-.%<*JL8-MH5[#!" $DI%(N@ 2, 
@ ,113X:7<_@V@FN;(X8E.A6"$:$)NMS.+/Z21!:A$K, 
@\%.,I5M3C &$;ERZYWOP\LP55:J]6VV8T),3BR&96OT 
@(E):">.D+,58,",V.8I2:!,J-7:'PV(0;@8[;DZ'!%X 
@0"(Q/*49+/>WQBU:1F%>BXG>I7:'3=05%\54;6:48D( 
@U][.^#J=2IRPE%KG"%)5"57BB0K_[9K 5W-^G$S7O:X 
@@3)X1 6G^'J%&!JA;3+-4/GAGW*43W#&#L(S>TR1@,0 
@U+?R;>61(=%\/B<J/ITT4G I2;?IGN<ZY;GQ,JD6\TP 
@6!(AO&NR(&K>N=-\-5Z3"PNBGF=X;>.Z9PG2M\\$1]( 
@Z;B*$ \K*:6\UEW^9VE)[Z<\/#UWM-#N$ =_ZA$4EFD 
@_5'>(E?8248&.6L[0\]^ZKX3V,H&_<Z[=5(!N\.;OC@ 
@I10$NRH^%&M@@(QD\4GU65(I0#,NHS"VPVDJ?'QE5@L 
@>QF$]C^MB:W0H=!8;S.[5*#&#]$G_-L/MC4@^<FLXA\ 
@T7B!$W]=F+0O V1],YOC1.2X*FG^_7BO4\?ES#9R5@D 
@H@,OX4MCH!_,C?(_%+KU#!1A?WYWD-PR#NCQ;.G(B<, 
@-B!#QG5\16E%>O09<AK-0J4J.?>V[0)G9*%J.BWS6HT 
@(&;'@;;U9*,!L%+W[2.5/@*^ZQ>@K:OJL2F=+L.LA]\ 
@+<?05_D['10\87?)5<PD:JY0'*=Y0\N,HVD?<F!-/<P 
@>H'R,.6C8@FF+))-V=>)2:B?;(48@7P2B9]'?C9 DO$ 
@GHS$ E U/W)(V:;L^K_[\#@\4@@--%C)3^ +N54E80( 
0#8EJB3&/@)1;G@M!KZ-T;P  
`pragma protect end_protected
