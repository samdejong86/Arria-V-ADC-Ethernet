// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
feP6IOiriiMOjRBiD/zKGseGwlSGoBh8aOZuWr22e6wR0vzs0lDe8FZfba7Oo5JxU7OLKax5JxLu
ezDHl+135YopVXdCeJLxbXqFrNgLpKkMWcOpACYfARQN4YRqc+9ZvKJ5HtYVabFxzQ+7HQpMUZLe
Vx0OLPzrGa0L/CfwPYqpR22cEQd+Sksw9jahlZDl+JGiR8diWwtefIFC+HXZnf6IqEKtqmexislC
H27I2xWIwzyi3nv92ri06HeTB7jK9GrljoZFL0PIcleVDPmofwESc3FjYN9eZFASuNdyeCishKgs
UXc19+zstYtjth3QsuX3w18T68hjAx1L4U76VA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5104)
cNnhdo92IVVM8Wd7LEMA7srVtQw5eZxJlpqUb+IszQKd1FZhSeCOsvvS7Z9s2ssx8rng7gUtU8MR
VINeI9bHj9eDfU9Uefc3lBFj9u4UjbDgkM88ujAoPnqpzWIX81kPXN16aPBZXssVmYyE5Kj9Ibc8
F1OHw5F+S9JuhWGrbYTkYSBGyfhCtXsNG5HyBhjjo8NfN4vJfQ4zcYQXCrUPaK2hk9q2RXP/+poW
XMb2PdpMbt/OXrizacJAPbZdQzSg65T00+53k6FXzcc0MeeREYFcIM5bEHqBGXhzSOqdYhwLD9yV
919BRePFCLOpNSIeVMUwQf9PqzmCpTJRYbcfKb1W6DDJSipPCL8ignROxz+hrLq5xXXYJfwGnc5V
ECl6W11pFsyaHx+TVdZLPOiXX+uBzYpNsjC1+DsV4fhZmLOwEsip3YV3eNr/HH5kUWT8Qwic4D7b
guONZhrk4pfNQoPkRTPLfSr1u7lonMz1OsDQBPR1V6OjrpI49BnD9u24CHpmHPrMr326rR5up3cL
jS6OZt6snU7xscPFKTDvWER0m75xbauDCLPyQMVD1TJ6bXXTHbXusUlI5a9Diix5b0ZcHEYSIQ8a
l6/jDnMy5d78Oa04SRJdQ+NFUYADZNuiKvhT5NEBd71TybP0so6SQWqYHKgquY6REmAQsXDaOL6J
PoMhrCG7qBESfOZFr/toSh/kB1v/NCuzuYLynQZ5DG/upPnYKIxB0NwQDMilYD6wEEMoUQ55wDfM
7drhK3dAQRWzyCe7y6fut00NWABFAgJq8vp7KDRL8uvgbQZBIF5CxHGoyjNzD9yuptFMfClk/KFE
+TsHxYVYod0FVpOewnVkO07hBpaXTzpZWD0HJZubx4kLFl4gJpcWVToorPKZCNqP4Pskm/hTgqv/
9RpsJHjRWR0+QxcrYVBjMLsiDPLHITMtkGVJeSjMs3RMkYor+t7twIv1DtjOZ+cWl47MoGyYh6CI
yfcvVHqK2wZwITrkjGRSBzJBsDjTdxFiaKNRiN38GkZ/8jxT0Rp0NsFo0ra3bcf7vghEg0/sMKn6
DTFe8KxMT2UXWel7RZcTjFWZX4xP6kvBj8a3CxvGFcUJXG/7Z+1PXw1Y6o5KhSHGabK667jb7tgw
dSdOgR7fSQjOz7MJ/RRdEddRLLFYsSJlNP4g0JVXrV1nUtryG5EgHZLP2gtYlCgtHFdh6OVSCX2b
YNl8PuTjfegeJ25nO4yeq64fuovHhHz5hXqQwqAsz+u/Xo0bQhQW5pt9s2tBP64UOTUW6okbZQ7Z
L3T8uUCmuTvYUShJm3X0UZnLqoTRMhVcgZS7KLFq8jiAqx5NnHN8thE6dqFgwtozOgFbAFsRgjhy
7XGHWd+j7s8hp02+RO5eRr5dWvi8+INz6s8xgMqhlwre9tUSHclro45Hb6YmL5BHirULNp4nFNTp
i1exlx5RALWt1CuSYFBHeRNKR3KC5b2HHgTk5N14ig4CiPDw1oGqQsp30MG3R+3DOlnmc5ojV5+D
DHiL/Uwi7n2ZgvMwWAFzThvqpy5JE9VG0TTyJaHVodaz2HZ38wiv6b34b+wX6R9wuo6A0fzs13II
uKQsGpud9MLu1ngSDLE3JNxhaUKTOwY4V6yHpNqKcYHVJv0IL4Zfca6CFQEMT/ITwwcOmsBoMW+4
yigAzOs0KeuTHWjQyAk460LGep6PQZqxoaJwv8V72Uq6m8CahfG5M9ZaFgacQ5a/BETfZ+BgSKbh
tU1uGukVXqZBSPedCz8HW4rpkFmQAoYKeB/ynTQLcu4E/Y11dyvN4EhNBBNq9gQ4EsBLz3lJbkJs
aS/QNKv4E0dmtxbbv8s2LzAQCKxin0VU9M7616JVaYDinfGW0PrRwX+UeCCMT5TGJM/zXnmATcXp
UcByJop3crx6L8OpQRaj3Pt/4b2CrY3TVOpzj+qsWpkcASytIy++uypmfJ9w5fUoPVFUqWtt2Pjo
gm7Q9GjN0vi3KQe5Yidy60j2BRMPCoaMZWxfS+Xfo270qj2sUknWP0lqb8N184PM0UrI4IkOrY8a
x2A4WLQck5DDKchi9TXyTBit0mt89onON1uH37k02cDQ3K0M/gX14FOpUKArqzZrrCEZvkCtVcqR
OAkhFQp75/oH9Lof8BABClgFY6dxuaTYOkfUYsDganWfzg8V+hOYPB5ftPd1wbI0xuQ7RVH2s6CG
mBMRx6dJTG0qhdu1ioL+WCf4boK11rQTL+RWY5ysnDlUb1XKWojzO90ZKFIiB6GuDl2D2mecEDWx
x9WROuLZhe+lK9hJtcmHMWqkpmR4P4P3kOm0wxbgG19Epm1fabc+8gWk63j0SmlLgngglgRKQxiT
8DGGRypEfNMI1oC3qSEml105z4wWyZiXqnN4wzALOCPwarMn2OTFP8tMoLzVinxCfTTxzxlWbsqR
Zs4vVDFDAXhUx98YjatxH5FHhslMRb7KXmIbhJQSGEp529U768qNVlBDJgFLFMx6fKWEbqXk7vGZ
NGmB5v98gFUTgtI+3cSARKlv1zNdSrPjHxY5IC0n4vZrJITlKUwAQ1kVdcCjOCoijfxqEhFb24ES
iidZQ/IImh8YcLvx8siSDzrvy6vkrw0dCvOq9yYEvagS6sSwR83sx8i9cXFsGAiYjAUjt/CxBkrz
5uqClsv2AbKpN9SzanIhosx8HYj58mVd8KggKxj+SoKUnZ0Com3jrZKNJU1nMyKO5oax2GQ9XOgI
R5PHZsZnuXd750nlmUDb4PwYzfzU+pZBu1rbiZdQPpuFEirMEgghXoY0jw2MPkCFA41IyYvTvnnP
Jdp6QYnUktgUiwWDZlvQ5ZYp0imqS6fIj6miShD+1hyxfLa42eEAJSrEg44JNDLdbEleytBaO9wG
JPmd+H6Dfg6eug2vwcHUdruv1ipJKlZcuwCtkBMtRZFVP6MMoqyWm6+0ihMmGHruH2qpPxbpWf4m
ooUBpnfRXxWRdjNW3B7aLdNEu3MKUGFXK0YZ9Vfv3Gk9VY1KP2IIJNse/cmyM4/4aovMBEk4LY8k
DTG+9UsO7EGHvWUB/lmi3wkGB33/wbdOqPTVArl+OPRUggL9mX0XoSlYuev4WSrWsbb0O6hFKpPn
c7VQEYZpKeE0EPgZBYq+OKmonyjf7IgpHpaG2/A+uJswr1wVAFIuaeEU8JZj8UhURQOx9bAuAILa
0k9tRJCS95V0MnYbQT3+0w+g5G6hiMZCxjBZXn0OwyLDYmNhwENf+A4fwtZEzmAkEUQ7aeDwHvDj
IYSt6XDIK7QdFVFz5fQWVcYB8Q+Xa7xnf62D+DdelHudJZ7c2u3s6j6+1Q53rkb5FB060v4261pU
6OQwWFA0P37N4AfG21MBuLPrFoG8sA9HykYYQda73Fuxxr48gouO3H0eUHJHsibmfchPNBPjIAGG
z9dOWuxXrnv1jtwFGxls6JmFWlEhcu2bc+9X02ONSJGwEEtrLk42Rv6arXTi+SIythIqdN95h+wn
6qifqZmJH5oPz7H1PZBA1bHcW0kbZDhWRb4NhuM9nqPiOCt7qdqjcKZ1w6dCZPdy0uI3P60ur0+N
5lcpVGpYrDvF8VAHyuwRYD0D0RBeXFYwp/swB7gJaW2523DaiGbOVk1fkcZDSqb/Ij+Ixc1qC1Kx
0JfvyMBZz7X4/58k4uNLmyi1rnGFktiT88YyodK3f9pwZ9f9jXwNVw5WcMaQds7OO7EU/X/vQHTB
mrJAcDf+3tRH0dpFm+uat+NltprXMlDDkEHb87i8Z8Z0nG1wq8SNUtyoxoh4pWH6sA5LAnlFACcv
WSn1MtlWC42bLohLHE1TpC23bjofMN+KnZVPI8i1EXWy3buKyN2kOnCPXMJwtfX76TIaJnBl3b4b
lIL17bFh1gIMF01Ve9E5lIMGVrIfs2gyYKyMZ4geUpVhnWdD4dyGEH7TwupU1gIBzqIbKc9yXLzw
xZLgIINrMaW2pbV+Hgnank+Iu6CnEaQ+UNWSD1z80jd8yfp6W0Pxp3BZvBNtftEvgwzTS1E59Yr4
vB3x4SZ1Hw7tpuykKhknzamiB+KH/NwCkb0sgf6LS32SXNjFYyGisnQF3J/XNh8UVzeMhsrtb3o6
1NaiaQdSfIrVGc4Y1Ca6OWx9qsPu78ugY3MDAXU2ljwM0W/YD2wf6EbVfCqhJHcmfPnRnXVwkt6N
16JuKIpgqfR+nOa95WLh8xrGTH7swHe1CPGVA9SyHu8XdfQj7zJMW/oCNS85Bluu9kuvOM440qY7
q/W8FU+nbXPMReDfjy+Mrc5rpuk1l/KTaiIOvarBScVXowi4TjXqaB6Njhr9DXaTjfX8t4DTKea5
+FWIcB5qOmNqkjAkbooBnR4wCbqtrlKQpJKaFm8SpEedLcIxBGObs6zDqaSa9y55knO7Vc7OtJr8
Cqehjaj9qfHr+d92IhDW70djNTZFd96rj6iZFHr53xTHz0TTb122pnU9G6MDu7VzsQZGqMXBqseh
+6ovlgN5XDzFOveqeOuj6hLZ4Sien+1Zn/DKJZF1YIQO2J93uUu6rEhUSSg7GMUUkDvR5ayKj8c2
GnUjpsJ8kZw2wGBMMLbTEmL3mK+C18GJXJuifmjCeXylBFmNEq51jI1E24kkRaGDzHHW1LSrS8fL
x+7KrNQkYZYCuPSIzRDJV11Nmrd7KfLBJz1bRqI4/wRmguhd+PspLJ5MBBb9q/zJOj/fmAyFb1an
AFah1V9iX6GhlsWQPXbVpj5vRLPsrNltqjJY5avWdJcOIHsS6Sez7Riz9lKDbS4tg9nFm9iJ6/ys
qcff0JsOF7bBK5oeBPNmcVGjdxCuwEOvPQDv3l6Xx2ZvjnI9CqvED7nK7RhJhlaMNBrRippz8eUj
7XTb2vS8wMicw+bhf5Ck6ytlcEqOEJAnjvHI3uxCNRc7xV5/ZUp7EKkMtFW2PbWO2h5ovCrCKcXm
TxQcPZeKdDTXBjjySU86Vs1yTMX+sOCtWGYZa7HHMlancRaR71H0fDCRDdg0irm8vmfDrEKeufH0
IHwCWpplWkh4sv4KXeHgydMkS+4fdbfu/CoFYpvcYOqoEolSCEC7gwjRgADZmyze6Eaf6YWeRaRI
ZSgYDqF31iQTLa1MzY7aGoAce0PJaBzHDnuNmfBIiOREJcytdv9gTp7Jo+WhDClIhhiL1TLAqlx/
2GPIFcM3SnYE0zgQibUAuewMQS2/6nJ+JYC3yC6vXqBa/tZqgD1pZgRAUQvysxyswk/fxGtb51R3
40+nts3C8LaYuTJfXrpb6iRn6mo7RTnyMKqcKfvhiH3fmni+C2anJtK7hDDh7yDyg/+a9van6n5B
LgxqlrLQcYOk8OgpTKuIungWJEAk1sFWbtmNBXG0kKs0Papd94a8mc0GJuOo4xAsmTiNsUkns8M6
AzxGdlQRdxRt9MEA0dgRarbxO/BqcuJtsHH+etot6/3XoCkcxs4CVOEc4m60U9e/170Nw3r+B5oJ
BElr5WUizAOmjr9B+vIVZsjY8Zpv+YAKCrNBTuCPvl6nD5ZpEZYLvw9CHC/fTc26rlkeI/j34kPj
Pi7V9PaZ18CMvu6A42/OSX2yBFiFs6XwLhUNxomAgmMbtUKZP/mzKAZd/Wak9114soH75BTblEnr
9AsB7aIb+BMnZAR3G+ilQqFylz5vYi4QnQPttds2xoDs48H7mkLVLdNsGReW2Z7E2rdpHyeqJFMV
yTtvRNDcTEl0hlNubJD/LhNVL6XZ28v3Jue1nu6sKBvdrs29XEXEwzkbNFkyIL6JL/wg//C4MmMv
Bi1oyB/9cQMooRXJj8bJr3mPcqQ2iEFpWFFUYmZnYNRAr0Qj4nIe4TL50T43X5cTSzNIjs+bAuFc
aJD6qY9mrfAfWIO9EZ+lPLZDMwL1WBUooQkj8uaWYqryfBj+A7AV8fDxGBUWRfqZGaMukMRA04sn
16LsVqR2pVM4NYA362EWvv17GES0ha8m5yJXnn11M/lkjOf5kR7jvy+ayGp5BGycV+zwhXwTFQUG
2VrkDlssZxW0T7ziZOnGZn694irV+ijQfxlzJ97/NozjJq134wVVEyl/SbwatOk1iqn1sXR/k6fA
FB64o5JTqeKxUmQXB07SLapvyCdnFgQjq0+ySQJSIaZPw8D5rZcG7V4qPhQU/QpvwPTNdZZ8rcFI
5yxqEJS1kvbIE7LMqQ+aLCxZpSasY2Xfzy4oCyDdp3rXPF8Q7qPZOUHhO7IJQrP7l/9CueQp7Cjn
QJPsrfOvhy+U8hAF5MvTQ/9Wv6JJNtml1nmnqZhAzJfghh5krP8+1eaL/jPry66nfxkJt7QjM+PU
/qbFkUC+xKfbPR/zcBsRnahWJVS8nMBzgj9BDCvTGdbFkiU552UF0Z4lkMlEGm+xPYHvULf5QFLF
Ay4sBfYddsXWXxBO3ZYm85ZZ36stjw/GeNDFqi+jE5bAD1847IUUQctfRH+Xito1eKhwk/adwCdA
WQfUB61k252ZguUgtC+aOP8A16fm2Ghp6Ya+59PZmlTjCVfkV0quWADYKJCewZLulNyuxJNQayGx
KT38wLgDWbiKgoxn7Wn+j0LDMFX6vfl/yD/iyXfhL9mwxpbJrkitTtDR0PL+4xk64ChGjrdU0rTc
DMelP3LJ3XT5Jz59Q+k/JH8B9r0IOXnT+dKrnsX9HHkAdMqN9I85BobSY9zPtHiTIMnlTP+wDdYL
MZyB+rAvScDh3Xo2Lb3ffW1bMFb0xLzqYp5me+2SZ6iRf3hciSvuA3PCSaNo2vxxSjwmucaty6hk
CsRfphAuhNN7rPhXLwEwnn2biYPek+nj++Yak1RZ8g==
`pragma protect end_protected
