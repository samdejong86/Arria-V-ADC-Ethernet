��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��N ˉjU���&�֑e��8d{X3]R,|�CbB��Sd˓��a�s���>D���7=ȭЈ���,WL�95��:��� F���Y�D�]c�0Te��Б��]��W�6tl��(~,�7r��5X���P��y�B֏?9�Yp���j�Iꘃ������i��͛�G�$��R9i��ᩙq�����J���}ҝ�h��]��0�*I���腏���E��8<ST �[:�R8��&#@�$����TKd�Ts�B�3�R�T����Jy������� ��H.���������^�����0��>�)�K���T=��{��|M]�"m�>����"��%7��yiW]I�F���0me��-Ә�Z�w6�O�(B�#�5`ò%���&�U^��[� �3�� �ލ3"��C/5@;�|$5�:�օ`+��2(�Ԛ��-��o)�� ߋ��|�@6Џ�4:��4<A���kU2w]�!*��n����"`���bX�����}��|~C�'s���`�|4>@�&_��uؒʉh 伦��A�X�P8`P���|���nQ+k�U��?B�O�A���I���*���4���K+5!�Y�Xr�ƄJ��M�5������j���hU���!\D$2�+�H�L�E��R�>1����%4�~�op��ú����D^��n�)T�][��c5A���=���B��d��氡�͖D��κ�߆��^$�Cȥ8��#I��?F�9��`��"��JZ5�<�� mY��
9��������J
��pH��:g��Y�!]�E�F1#��a-�?�R�_Ux�Dj����S�����7���?���x�ߌc��nK@�Sk]�Ki�6?�ۡ)ϣl����%-t���3�'�ko����Q��s�b2���k���"�y�bΘK���c�ܳg�"r�_����3c	A�N��o$� aF�]4�>�����}D+N3�/~D�����u�b���)l:�x�G��Hc�ϯ֑���i�=^*D�t�y�X)b�e��M$8��4h$(8p~q�w?Џ���V� �q����J: Ө���~�W�#�M���֛@P��LI0��d����:��(X�%SđF�C���t%o	�X��e�3�D��*�R�'$<�,�>�pM��ƂY�������e��*�E�����3m��V� �Ξ��{od���Y�{	�pnC�~��9�zv��
?�T�`˸(9p���.g�E��66C#�r�Ccj��o�NПi:h�+�~"7���������k[�����B�Y�ƧlM�Hi��I]y��P�aWu�`t���$�X�k����Uon=.��U=w ����0d�QJ>����ebB�6��X�mu8�y�1���m��2&{�����IP092̰�]��eM�+VD�Ear��%�Q�)���+YM�3�X���@�r���VH��rP�=�|��%�P4(��u4����ˬ��Wd����k)t�r��H^�PX�y��#?qg���{���	-�_����>���-woh��c�J;�[�N	�]�ӣ��<˾_{���P�P�7����g49�Ws�rz�\��V�H��#�L�]���$��^���C�2"uqF���V0�`/H��H�����a�Y����d�s��!0�zQ��t�����\�p���U]p����\%E�-p�"��My�sz�.���Ku��/��lj`	t�
��3�F�EÄ�xe��z���M|m�[��ZLXF���W=U�ÏS��ì�f���q?�oHMM��5��"�-*X�])�`�ÿ����[V���dG%�4�c�-�쳃F��(��mx`1�I�F��d8��Ŗ�!QZ��y鉡Z'��S�ş�UO��Ho�C
�_������o����4Md_�,��e��p�����������t!_oV��}�w�����a,�`(��"m�&m�v2����b<�>^���`��3aY�A�Z<Ӵ���#���+��n�������Ϥ���G0Ϣ�v���`<�2m%Ԯ擰X��-KҪbFO�Tc��?2u�ݲ�E[��c��b����H
��QV����N�SVM�JE��ڤ�w�]N��ek�=�!�1�/gQ���ʩ4��zȏ��ÖU[�>�ri��g��t���'ZQ�̺"�cD�\N�E�F�Pf0d#��5P���@�OQ��8+��K�J�]�^;�ɘ�Mlp���C#*sG�4|�|R-MV�\���9=[�,Y�bRm�3��\��&�)�RMCX��S?�Q�������>����o��>��4�����|��2G2�T�p�B���$!�m�����\&����_����ܐU�wB����}v������Jl,�l�D�挥��nb��]�={�}J �;��۲'�1ky-�m�0}c+�A)�o�S������ƹU������H/�S�J0)��?s���r?�S=&��] ��3b-�SPYut^m��a�]�/l��^�]�,��w�q�ip�P�do�ţ�(;�!Z!�m���o|گK�w��z�E�%	-�Q�a@�Si�1���S-�j2S���#���{BЬ�����yD(���fC7���P�\^���"�<dB+,��e7&N��� �ԢP��8�0����9,��;v�e& A�M�i{����Lj�X����]��e/Ki����F02������"Pʶ��)劒�W�:�x�;��D�%�)��C�P���`�ax����8�����v߽yyu3��fP.S�}��֣���� i�5K��Q����0a?BD�2��C�h����/���B�!�ے!~�/�zs���Ҿ�W�C�ڇ��ةs���Z�p#�xV�J 裚���3\����8
�`�~������l��~�]��]l����+�~HX�m+u+�����^��+���y�7�~K:5�^���V��ᭋ���Z�Ă���T�IY�������]����al�9!p5��$�FWN�
�a����4Eo'�.�6��iC_?�|�NPeA��R�����]#���O�������X2�)&ٳ�*d��|(V9�p7'JN}e���2�-���I�TJ�glYKv�ba��fv�ʲ�󥡑��{����=#b�8*�pL�"�E�����!O!����r1�^(�1q�	�>��1�3�X}2t��Ӄ��Ct���'��������i6�3F�f�0Xn8j����"���T_F[�}��r�����Y��	>�Lk�{z:�,}���@��k;˦ *��ߣ������h����(\!_������\�[&b��uG��H��!#�����lH�Q}Ҷ�#j�4�-�ŸؾճGx[� ^ԕz֞07%Gi�Z
��U{�3.��ᓕ��*���'�<׍e�I�j�۝� .�����Ye�����n���"
"z?>d�︥Bf]��%�ߺ��)н22_�S&}�]����
|;pFs7w"�L1�"�u�%��L�I���a�L,PbS'DF+˴��֙7 �oJ�B��%���!�?�c�q
{e�M܈���"RS��8���専��k�Dn�y�F�ǋ%߰#P�OH��p2W��Bwb�� 4:��{�I�7��cA|a��f��[{��(��������jLZߝN���0|	��D�{�B��v�< ��
r1�����(?��a��������k ��[BR�[l�O�yL�.��:��U�ɢ�}(<ZZ,��_�Y���]W�h�YC��X�`�?8�>(r`��7H���*�'��)��.�_-1h<�Ą�Ph�/A�;qC��2�̎aXYHo�P�
�:���Fzy��+�N��:� ������J���s�u]�.���w�>����3��p�Գ��>�Ja�Td`q>�#��~� �M**>�DTd����I��t7H_B���@"���X��u����CWJ�> 4���'|�>��0+��ӻ��|����e*Jh��?��ҁ� rԗ����T1c�*� bo���Z�`�g�>b�¼O emi� ����I]�E�4�Q�`������Dו�yw���A���|�/�R�F�%H���t)4�M@�|l�T��������n]6JQt�p0�wOuoxs�����憉4�� 0�*��(ޣ��b����n����ح[ME