// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
pqkOwfqJA1ClV/pIiQhl7C/PHmOSTyokF2OtcjYFwCzCohdfg9Q9Bk2SQluAaHPMsvmCRFx+ItrL
e05TJvVhvJtLARafXPHqRGw3kQcDFGCwcLF7VNAbNpe05LQpMt87f8WfrdraKvwrz2PdCGKkEVpz
zrmsr9CLpc3YBNoD1Wj5LjUTQ5XFYr+HWKWIYQaUoy22Ncp6JGfv0wcep4plmgjvQ8Gyq8UXgJId
AXjZ/s5aKwTRgjWDMqMVSTbbrby+6Kt1kgiDOacCbVynyx5OxemcD3A2Ou+pwL3HUFPYnsn8fPcs
GfSBKV4FuPhML1UB24cl2jvuaJ/BJ7P5G8kcUQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5600)
28NKPaYeoiFritdUO+kzOrwo9YeYFSEzyeQLGTxh3iubUYp8XWT7IVBDwIYxOCrf+Se9pACoCbpH
P0FbKL/3DMW5E/zY2/380X9184ogRkuMEyrv/T23KCn585HThzv/grHkW5YbzOrgAY77OF2tY1bE
KnIiZruKRDEMPMM++iUim3LMxuPMpdXEyzOXxeHRm4CZANOlTdm5kst0vPBGBMKYarNv4PLRecKc
PB7G5H9yhHP0bgBVoHjD/g+iO5tz9ft1LxFNAPTc7DICogeaxB7hGUAliKVQDuUP1J5/CNQjLuvE
8XXjl4+Xvd9/2R7hOObnQvlJIuobwiffi6xSfGos/7fHVlGtwuBF9IU4BKT+8FfWHe7nXH16yDUE
D+xxi+a+F9H2HoMgh8YXBYfNPRD5eosdqqDHTULXL3QjIbyNXzwnxPfIx0EOh7r0m/Q1cwZZU5zb
Ozz7YwUdgkjdW7wMAxgoDZNXWJze3MHVCDnZd6cGxoMQRCxEEdDzPqe6awQTC0ELeco83zVRS1uL
hnDQYUwSsSkhN5RhnW1Q7EQARHPFB1eL6dZcqNC5ti0yZ2kLTkjRuNTw2IQPwxGMWvIvW1oIagL9
IPa6/1UfGZXjr4XRNO2zsez74TrNPjc0ZCjY08aeJrHxwhtvaESVVChQMqS0592tEojAb8pJhEIH
Ui26EL7VfsTDL2Thiaj83KrrXOKRlXhMAOkBk+70qu4SLy8mEz6/VdbNFKHb8jP9Sx1sMDEdncRK
gWuemEC5iUFSBrm3CToeZw0l1c8gqamdS/xn8bXjxcK0OtXPrtiA3Bu+zjhcQ1dcnSyC0Mh1D0tL
7pglZJAm9O2pRubI7Ji7q2uMFw8+anHTt9GvUD2w/0pEpEAL5hXguoYvzC1632sE5U1xUvFk4/gH
/quoVp7ou5KDSY8kvYg/xg1zvAh8lBkmtw2355vqdvJhI0Dp7pKb+85clPaLWphfY5xyeMKO1w+6
LW8QdS8QJU5Fp3m37UO3IP/vmYJfgRAIDpXfqk31j4TorBEfmGZ91h6QWsPJXXRzfYGJeugPlQik
pqHnqI4BI3mPNdHEkoYc2ax4cPRlt7ZWsnHLK6/8SA7cFyKeS3MvhIwP+PVDDDuDkCXJjNT4w4jv
v4qZH1HF1EOM+ChmLRJDLoEHwKT7W+NgxikUKkK4BvL5xsKcclumAwGMBTJzy6haSIR+2BhcKoV5
pcRCWlnU7Fd+Kel7Q9UoJRxRWANmdyR40bHnuntbe/HTmTV7JZ2AJ65NlGstmM/0KrnrP4KzMRp5
WyA4Nv9whREzgV+e5/0HSwdyJSOj9K/Yg847Mklf3dXNZmDQdyDLFk3u+0K60PS+Rbk54ROO0PC5
O5M1oSFYb1VbOeKoCVn7XwE5KOa0d09C15pzOOxYxX1GlwwRsSIR/nrlw0N5wheqve8a4y6T3wdU
RGzPRQadRRm1sHrBh0xU9LmUrZItYptG6QSb65s1aDwdSVh+yniXGvPWJq8WHXzee3Q+tkkvk4hq
3A4kZFycUjlVa+gvYoRndDsaTjAVlHn8yfGXBFnn+XKksnNVcaoxQOqT+O3zBVKLA4b9CCIRam3Z
cX4T5fATEqe8CVxIHSDhcdBmjjSzw1qRXiLr7PUeLiGYY+FGEZVbv7EJxQfO6i9lrEXUgDdgc0Ke
PEFp85+aagT1pzi1ESZfOasAV7Gxz4GL0P8XdRxnxbEcbyaziYzCDyCuhan6tXBsfUGF2jYMPHg4
RrrCApw54ep4hX0dLluwI3izi0H+g7UKmYw1kyq2D/HcdhR4f9v00I3YiAEG4GkQ2GsHlVo8TwyG
pHmqAFeM9+Vwu7bCU3qlr/c7aC+AwzjPuA1ArC+RiEEJj+gtaDAm3Be+FTCBMFVPDqR7x8Y7zCON
22mGBpRWhqZM4OIf1VLCZyEFMkq5wdBAhmk3RKMnuK42N9Y5L6UcATdSmtF/03b2w/Cwu7yN+mXo
zjDImuqa3SUfDYG/SohB+az5JSIJEwVSMHofBlmcRMSM2Uk99/RDF96dZxx9qo0O5jhTZiGWJICs
D+OZ3fCB6FVMVk4BOjda0RKGfrclEpAWuQxDEotDnbBUS3gsKi4RjEvEQocH1DR1UxSU9VweLS/8
/KwBXzDMGhxy0sRvvmivko2pmsa95+sWoT4zFObHaImvufj8TW3XY7FDqZ1UZh8OtNPh5rZJqCNc
ungvUzUvdgs7PItXNcZOqLl7z1CsoE0gwhUUXY4eJ5YVtqE5SAgNh3wFTMK4oC1JhTX9zWQTI36v
BhBAwf9YoivdOltyEl4v2TxR6QV5kduhDurJtPB70P5BZoxVAYrZ2lzv3Qfy6GjzFOCLi5ZsKgfo
/ZYzOkz2Aqtrfr/guxD8OP5Vf/+n0tDu5aUNc9BiDY/dFveuX39yqv4f82MuHU+PaVSo4X9kzMbQ
zaLw7FwuP/Mza1HIiZdlbF+nUFiY3oaEq4dFX+c3ANao2PgxAs8hdRcEMGOb5LURL3bZ8jYJqY03
rNj5KszjO0Tt6gwNw7QFoS5/pEOSNu6JJ3WPbB5x2izO5/R3cFjtDM7r8zO4iSIUR0+txMWHEkNw
S/9Ca25+ThqL2undWAmoDZBNdbXUTW6XCu72ePE5GAaLTV9bPvhwExD6T3r7ny7mNdQtCux4bMMH
RC87bLiklXuHZ55nIRH/BlClU5CCZNzc+eT2xYZHyQMnVlHECQ6m46/wav2NOfaxQRuaCEd/jp5e
vhtAGZM3aBFZnSqEAgo5416FTlyIIRyB2soFon+/F6wQGCWPTfDJ/K5p93pcyQmVFWRaNs2fHaPp
pSupjHYjt+Y3eZbFPnBV/xGyqCzaOWfKpnZJHOiN8UmXVKmS35pmy88+UIgDJrMsi5GRk+iD+RdX
yO5YbLRoD8mA1efCYTcGGE53rBI7n7iFp6TNUggyylpyt6cv4vYYJarQLjvjkwogblIuFRmTzrYC
gtZeOzkl8F/tnLAJ1B6++obTS3U0TGhpVEQsvkYz+0ZJVf1gFmcFwVvXYC6tyBKlc1UGDaYEFxZy
v/43x+1uZBpkESvWpfsRRkxThY+RrK1kChqUCvHbVhQJ/uesMvFUgoL/murGvWBLNjKoScFnAuxC
Ibm/VmMFDHWNw4JydABVQoB7C6nPChVxtzSAjXAN0J8FXnLx07GjtOyQAl5nLEnEwyL47qlxD5h1
+kKkgXxBh8G7diH9mFNLHMxI27tpJPciEUFp3TGgwp6WF6Rz9YXxuwEVcgn3XseD8uJ7h153uqzP
pdQivzKvY4zGB3Q+II2CQ/THHYUKhox5W0nBbVG9y4bjg24tvRxvC1DM3vze2UFPEYGvEyq/TiAv
+i0zV23gDfaUTARUBccfHT9mVEZHpLMtp3j1SKAd/11DVWdZmrvtnJHXeN8lYQcX1btmh5bPkeUB
xphRnDsuP9SLq0wayUf2j8nUd8z0PJgx1vTEDJbXQH6+VfMEGT40QDEIEVp3hFgkX6iv7gS+qlAm
RrlLEDMrPxw83Pc5q9QFLn2855NSfSSooY0Vpv9tJ/xX2bDrK7MP98rQVh2xIS7DpMtiii3oifrT
hxH/+nSMl6XCZEomUPliSPm4h6xjTBaFvNybUC73AeKbqOYYTDYCga86RBgDO1EUOqAajYT8jVek
0AcK8IGM9JgPnbG/JaCkKg1d7u4JDyaj0k+aFGkAAVcOHbxpiP2pnsviVte/hz+eX3cSrNgZTBYr
BuXiLpRMe9sNc7K1bQdkXAhLHuXiK50ZD8tmx48Lp3jY1Ggjboe49OQEcRX+pBTT51o2gdO4XjUs
CnjL2Imc04F5FObhtb27y4pisMtyUh04QroPLydRoODoBvA3IRCf412f6w4Y72SN25Ihl9yQa/V9
mMD3MTFpZkcqlYjg1Srb/kn3lx2u+Jhmgkt7gacPlPSvj9SVquP0R7+9pRgKsu0pbfxKkL6pcXAm
B3+E7CHKJY5aUKS/4Fo10d6j6tYCSDFbYg2cuLBAgbpE5/rVl8/VAv5rfeIaHzrub06t1XZe+k6v
zGpUoDC1xh/FTtZ7CdMfw+xXQHebzmkgry1u7RaUXw+wFN5J9VYozXMFWJy097syrV4KLzNvs/WR
xsHXNVxs1ohOYPz5WQh6H/T9VL8CwfFPtxyyKTQfeRdCW+bjAYIsUNUicPCHI9br30IL/O9lgtOP
kzeM7ULmdrcYjmngopTg8RGmJKIfsZf2ezWzdRAOv4EJcgyWh+tp1Mjlen0OmHFIyeTyQ5NauCSo
NC1AEJbHBrWjRoCKXJ69xKsz1K2OL1BwrrQ1Gp29Uu4N6RNEs31zKDRbQaoDP1oUSOHnUvJxnEZF
ACHdo6onzL9BRxhwCYvicbwMKVSphs5Ryy+dxqfzrZsEC10bBDYbMN/6Bt+EliqzxCeJ1MzWNijb
LKALVN7+1RifnDevMUossgnHWsF5IlrPeLO3C4GAOLk1rNuyz3NkJOAjI65pZzCGELxippX4tN6u
vfTi5KVb1siSQlyDTdoDi/U2WOOrvIbd7w/T+AsffhI9Vq4j4KnxJHm54HxOcwsP56wX4elELlrH
c5lLCnQpHMSFbGbLn3btwQIDLNUXydXCR0sRPOzmYBAnblzTWJz4TT5+vEj/a0wJJcB+k4jHQBVt
pPtZIpZogLtSfT3xCWYRyKfxeILVz7xTahl80GEOtz+zwb1+N/PuRD3osVP5ZO0WViQu2ZMXvFy0
drr2ZFVWyw9/XwSjQzmKn3jZQHlxzHl835CsAFXcC/jfj0kw9cea5fW9iXa7k6LgCRjvaO5WotQY
wm+tOKRg2Q/qMybKlcWmHu6q20GqDwpRdKCQli+eOXTx1sE2sE9XPpcFsnNE1uyXGpQUwjtsYmWb
VsnOcJbjl66y0WYs6SZbIzSWkSe+zpMk32BYHfA4inzlsuCx6462216l18kIAfGQJf6O5kbraio1
upKM6aQ829x7LPe6SmxS52q5lIv1KVsDSPlnqHhD7Or4AJhb5Uzk0zB5cJ2nBY5hBfRjr931OnaE
fNtY3LiKc9bGTakEW/PgLq5LVyEp2w2fwGX1F/eVzkUOYCox6q0Ip62Lf8DCJROom2nnzutvvVj7
vbJobfXwxBXCk3IP1X4TYjH7ck7c1A02z7D3WCabp2LtD1YsPkV/4gK43Vh2RchHqlyEurkh9iL7
rFBuDP7eUnbeuXgRrmC5RdEJLF+IqXAmDfljwwr9gO4aQlJ92cjqzhhwvVKhFDhVPQGw9ISXhzp6
RZPKQgH8v6B7pZaAiTgryzfDo6KX0cmdsBJOwOyOexp2emfLRQVTC3SzrTd892w6J8j7zn78C7Gh
5IkQazktdNom8YQXFAwXqkiVNmnlrA1fi+CYG7FZzVeU8yYxiVaJ8Sr4zi0pUHx2gmP2BAA7ZoiD
weKCeubPtWAU5F0k8HTdkeMVPUzLEl/td5qKO0Sf+/+l+7sUVHZoI6bfjLNS/ReYoC9ARZg65tbF
T4BLyZ9pcPVRSBU2W73G7o0mHA/onmcgebPv2sm+mNLECtZSi48yGcjOPLkYMdiG1kFdz7g5T4jr
QANnz3kMPGsHGA9B63Mtn3whFmhaEhNhr3afEQsDysTGbnIDUCE8CZYNqutW1u7m+jQLiuCLXeZK
qHItA/OKtT43ejBaGB8bQEcbl6AFE5eQtlqMqMR47nP8bR83DhgERhEX21YbjYchjWBgW8GjaGY2
VEt6+ptDd3TJmKKQMg6KGyl4sh/4W9+a2NvvPQDOayqUdcGq2aiUzMLj9+FMZIPJSvdwD1eUI7nM
1V+/zY8YU/LvWXlnm8rvUYKcfpekaeJcbg3Um+23m9KIbV5cFHkYg6/MIVp5iKJmmeTr7gC/h1Gt
0u5f1U246sYFvroO0u+miJBUC6eLEyuCk/fkQ3xyqRIy42iRJTAo0Ll+sD6RKWOq+IoAwD4/5qbQ
3lL/LztTWaMbRUEKCqK28bm5bCK4zyjfxP7b0irulH3mUcLQ3iLdHkXKtcyZA2SBRc5gRJElfqi6
wcHac6gCKD1bRDbQMb8N4gyGMPdjNKbPhCoHaOYScMCsAjze4jBTaINEZ5Qz47yY0H7YOraJh0bI
SwyU5+waKjreQWKoy5+HkXFdf1aIPrxvK+FkG43EgdVV8iHpvNBXGBr2lCEI4TCaq3DmLmB/zVZe
pFHxU4MDXUIpODSy9NiolQy5q8v2kwvZK8PM1wnxKsIFJl/POz36Iqp4cbKbYajyKWRAfxJoDkDl
8jKU6PTTCmx52+VdOXG72pY7IJfy2L8rFlmGI68Bk5cuG4IDDX9Vr2wNiqKlZdvJZJrWPcyLtyM1
kBOoJ7ZRptXvxNkdWOSsV+VTim9iOPlMsu1Lp/syyJb3sjX2fz/ujU0sSSyWyFYFARyxuxPVzKYL
DFnjz2mG0ormp6HHPmPlGJhBMxphEDjWArfbj5KPy4t7d6pcu9aa6HZ/NM0NxH0i6m4pz4r/SEOB
rtp9C9MrM9IZ1TZ/oxfEyJf9f2DWsioqiDsGW+F3B4wuV8bEIIUy8xqFyNnpnE0hHT8BrEtov2T2
eb/N/lPwRZDRnMoL7ym1UNi7/5fhlikwyJbIjCeh6lpm51V/pK51Php6t0Xm5E5VtAFKx9jbjSom
ZcKzEdfpYOLebbX4fOh7ZOccrbPvWa1cKjr2sJ+bych/YUsEcflKbLxfx3cuvuWyb36UI7nnpnCJ
oRsLaCy7DdcI4Ex7oO31NuXUY2coWUBKU+lI1Z/WCNWOsSh18Hu5EFi0b7pSq02xuFEfcE13aS20
uPss01ZPCzAeNgYEgtv7pEenjg3zDAx320VKqJbPlwZFmJO0p8WTpI8sn9OhQB5u3RXXhZILsq8Y
UqGI4NG22/a3DfIli7tkTuto6BsL/EdJpsyS7x6TG2tpNWiGva8nSaSqgSW3GAlLewR+SruT2FCo
5pWdNYlZAdvYPeGQDMevwUik43bZHuORWkpo49SwbQKjlt/qhdT+0aDA56+985bcMWbNvGTAAMz9
wXYjTtya3kgHXNOiSlE7GcB5RjtomFq1C4RXsosOhL5q/4w3I5ZOeK1cXy6ELf+dWzuJmBauuKRQ
NrNqrxmEcKNjQ/KG23df3gW6r9l0AkJdjHNhS32EkKyhDBdJBhYUWVO+gw/rGNHdRF0RcW8P5wDa
PSq/oIrm2dzKYChRwU+ktVs8lsonB8zLMW4VGA5VxQHwIbFgEsWFyduzWZnBi4Q2qRbwEgzbP2WL
vfcPu1avBWGOi6vveizos5+VEyfDi573xcxCelb0+WPkNcPgjsGHrXgKvgle2BByEo3QHfSIgrAR
AouxuIXC7pEnwW6miLzr/IhcVRBo03egGOrO3/8oPjAwJH/5lShut/rkuVOgUEvM0fmgG8jx+o/b
J9Dpwp05/X0M3C4FmCjGqN6U3P5UqONdrGKuEwemzXt5/NCZ7wjfaw3Wcukscep1/3xaglkGcOF0
qGPFCl8BU+LHDYvCiP4=
`pragma protect end_protected
