// Nios_CPU_qsys_tb.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module Nios_CPU_qsys_tb (
	);

	wire         nios_cpu_qsys_inst_clk_bfm_clk_clk;                                     // Nios_CPU_qsys_inst_clk_bfm:clk -> [Nios_CPU_qsys_inst:clk_clk, Nios_CPU_qsys_inst_enet_pll_reset_bfm:clk, Nios_CPU_qsys_inst_merged_resets_in_reset_bfm:clk]
	wire         nios_cpu_qsys_inst_tse_mac_pcs_mac_rx_clock_connection_bfm_clk_clk;     // Nios_CPU_qsys_inst_tse_mac_pcs_mac_rx_clock_connection_bfm:clk -> Nios_CPU_qsys_inst:tse_mac_pcs_mac_rx_clock_connection_clk
	wire         nios_cpu_qsys_inst_tse_mac_pcs_mac_tx_clock_connection_bfm_clk_clk;     // Nios_CPU_qsys_inst_tse_mac_pcs_mac_tx_clock_connection_bfm:clk -> Nios_CPU_qsys_inst:tse_mac_pcs_mac_tx_clock_connection_clk
	wire   [7:0] nios_cpu_qsys_inst_adc_control_out_export;                              // Nios_CPU_qsys_inst:adc_control_out_export -> Nios_CPU_qsys_inst_adc_control_out_bfm:sig_export
	wire         nios_cpu_qsys_inst_enet_pll_locked_export;                              // Nios_CPU_qsys_inst:enet_pll_locked_export -> Nios_CPU_qsys_inst_enet_pll_locked_bfm:sig_export
	wire         nios_cpu_qsys_inst_lcd_external_rs;                                     // Nios_CPU_qsys_inst:lcd_external_RS -> Nios_CPU_qsys_inst_lcd_external_bfm:sig_RS
	wire   [7:0] nios_cpu_qsys_inst_lcd_external_data;                                   // [] -> [Nios_CPU_qsys_inst:lcd_external_data, Nios_CPU_qsys_inst_lcd_external_bfm:sig_data]
	wire         nios_cpu_qsys_inst_lcd_external_rw;                                     // Nios_CPU_qsys_inst:lcd_external_RW -> Nios_CPU_qsys_inst_lcd_external_bfm:sig_RW
	wire         nios_cpu_qsys_inst_lcd_external_e;                                      // Nios_CPU_qsys_inst:lcd_external_E -> Nios_CPU_qsys_inst_lcd_external_bfm:sig_E
	wire   [0:0] cfi_flash_atb_bridge_0_tcb_translator_out_tcm_chipselect_n_out;         // cfi_flash_atb_bridge_0_tcb_translator:tcm_chipselect_n_out -> cfi_flash_atb_bridge_0_tcb_translator_out_bfm:sig_tcm_chipselect_n_out
	wire  [26:0] cfi_flash_atb_bridge_0_tcb_translator_out_tcm_address_out;              // cfi_flash_atb_bridge_0_tcb_translator:tcm_address_out -> cfi_flash_atb_bridge_0_tcb_translator_out_bfm:sig_tcm_address_out
	wire  [15:0] cfi_flash_atb_bridge_0_tcb_translator_out_tcm_data_out;                 // [] -> [cfi_flash_atb_bridge_0_tcb_translator:tcm_data_out, cfi_flash_atb_bridge_0_tcb_translator_out_bfm:sig_tcm_data_out]
	wire   [0:0] cfi_flash_atb_bridge_0_tcb_translator_out_tcm_read_n_out;               // cfi_flash_atb_bridge_0_tcb_translator:tcm_read_n_out -> cfi_flash_atb_bridge_0_tcb_translator_out_bfm:sig_tcm_read_n_out
	wire   [0:0] cfi_flash_atb_bridge_0_tcb_translator_out_tcm_write_n_out;              // cfi_flash_atb_bridge_0_tcb_translator:tcm_write_n_out -> cfi_flash_atb_bridge_0_tcb_translator_out_bfm:sig_tcm_write_n_out
	wire  [15:0] nios_cpu_qsys_inst_samplenum_out_export;                                // Nios_CPU_qsys_inst:samplenum_out_export -> Nios_CPU_qsys_inst_samplenum_out_bfm:sig_export
	wire   [0:0] nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_bfm_conduit_mdio_in;     // Nios_CPU_qsys_inst_tse_mac_mac_mdio_connection_bfm:sig_mdio_in -> Nios_CPU_qsys_inst:tse_mac_mac_mdio_connection_mdio_in
	wire         nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdio_oen;                // Nios_CPU_qsys_inst:tse_mac_mac_mdio_connection_mdio_oen -> Nios_CPU_qsys_inst_tse_mac_mac_mdio_connection_bfm:sig_mdio_oen
	wire         nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdio_out;                // Nios_CPU_qsys_inst:tse_mac_mac_mdio_connection_mdio_out -> Nios_CPU_qsys_inst_tse_mac_mac_mdio_connection_bfm:sig_mdio_out
	wire         nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdc;                     // Nios_CPU_qsys_inst:tse_mac_mac_mdio_connection_mdc -> Nios_CPU_qsys_inst_tse_mac_mac_mdio_connection_bfm:sig_mdc
	wire         nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_tx_control;             // Nios_CPU_qsys_inst:tse_mac_mac_rgmii_connection_tx_control -> Nios_CPU_qsys_inst_tse_mac_mac_rgmii_connection_bfm:sig_tx_control
	wire   [0:0] nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_bfm_conduit_rx_control; // Nios_CPU_qsys_inst_tse_mac_mac_rgmii_connection_bfm:sig_rx_control -> Nios_CPU_qsys_inst:tse_mac_mac_rgmii_connection_rx_control
	wire   [3:0] nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_bfm_conduit_rgmii_in;   // Nios_CPU_qsys_inst_tse_mac_mac_rgmii_connection_bfm:sig_rgmii_in -> Nios_CPU_qsys_inst:tse_mac_mac_rgmii_connection_rgmii_in
	wire   [3:0] nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_rgmii_out;              // Nios_CPU_qsys_inst:tse_mac_mac_rgmii_connection_rgmii_out -> Nios_CPU_qsys_inst_tse_mac_mac_rgmii_connection_bfm:sig_rgmii_out
	wire         nios_cpu_qsys_inst_tse_mac_mac_status_connection_ena_10;                // Nios_CPU_qsys_inst:tse_mac_mac_status_connection_ena_10 -> Nios_CPU_qsys_inst_tse_mac_mac_status_connection_bfm:sig_ena_10
	wire         nios_cpu_qsys_inst_tse_mac_mac_status_connection_eth_mode;              // Nios_CPU_qsys_inst:tse_mac_mac_status_connection_eth_mode -> Nios_CPU_qsys_inst_tse_mac_mac_status_connection_bfm:sig_eth_mode
	wire   [0:0] nios_cpu_qsys_inst_tse_mac_mac_status_connection_bfm_conduit_set_1000;  // Nios_CPU_qsys_inst_tse_mac_mac_status_connection_bfm:sig_set_1000 -> Nios_CPU_qsys_inst:tse_mac_mac_status_connection_set_1000
	wire   [0:0] nios_cpu_qsys_inst_tse_mac_mac_status_connection_bfm_conduit_set_10;    // Nios_CPU_qsys_inst_tse_mac_mac_status_connection_bfm:sig_set_10 -> Nios_CPU_qsys_inst:tse_mac_mac_status_connection_set_10
	wire  [15:0] nios_cpu_qsys_inst_wavesample_in_bfm_conduit_export;                    // Nios_CPU_qsys_inst_wavesample_in_bfm:sig_export -> Nios_CPU_qsys_inst:wavesample_in_export
	wire   [0:0] nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out;     // Nios_CPU_qsys_inst:cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out -> cfi_flash_atb_bridge_0_tcb_translator:in_tcm_chipselect_n_out
	wire  [26:0] nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_address_out;          // Nios_CPU_qsys_inst:cfi_flash_atb_bridge_0_out_tcm_address_out -> cfi_flash_atb_bridge_0_tcb_translator:in_tcm_address_out
	wire  [15:0] nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_data_out;             // [] -> [Nios_CPU_qsys_inst:cfi_flash_atb_bridge_0_out_tcm_data_out, cfi_flash_atb_bridge_0_tcb_translator:in_tcm_data_out]
	wire   [0:0] nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_read_n_out;           // Nios_CPU_qsys_inst:cfi_flash_atb_bridge_0_out_tcm_read_n_out -> cfi_flash_atb_bridge_0_tcb_translator:in_tcm_read_n_out
	wire   [0:0] nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_write_n_out;          // Nios_CPU_qsys_inst:cfi_flash_atb_bridge_0_out_tcm_write_n_out -> cfi_flash_atb_bridge_0_tcb_translator:in_tcm_write_n_out
	wire         nios_cpu_qsys_inst_enet_pll_reset_bfm_reset_reset;                      // Nios_CPU_qsys_inst_enet_pll_reset_bfm:reset -> Nios_CPU_qsys_inst:enet_pll_reset_reset
	wire         nios_cpu_qsys_inst_merged_resets_in_reset_bfm_reset_reset;              // Nios_CPU_qsys_inst_merged_resets_in_reset_bfm:reset -> Nios_CPU_qsys_inst:merged_resets_in_reset_reset_n

	Nios_CPU_qsys nios_cpu_qsys_inst (
		.adc_control_out_export                          (nios_cpu_qsys_inst_adc_control_out_export),                              //                     adc_control_out.export
		.cfi_flash_atb_bridge_0_out_tcm_address_out      (nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_address_out),          //          cfi_flash_atb_bridge_0_out.tcm_address_out
		.cfi_flash_atb_bridge_0_out_tcm_read_n_out       (nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_read_n_out),           //                                    .tcm_read_n_out
		.cfi_flash_atb_bridge_0_out_tcm_write_n_out      (nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_write_n_out),          //                                    .tcm_write_n_out
		.cfi_flash_atb_bridge_0_out_tcm_data_out         (nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_data_out),             //                                    .tcm_data_out
		.cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out (nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out),     //                                    .tcm_chipselect_n_out
		.clk_clk                                         (nios_cpu_qsys_inst_clk_bfm_clk_clk),                                     //                                 clk.clk
		.enet_pll_locked_export                          (nios_cpu_qsys_inst_enet_pll_locked_export),                              //                     enet_pll_locked.export
		.enet_pll_outclk0_clk                            (),                                                                       //                    enet_pll_outclk0.clk
		.enet_pll_outclk1_clk                            (),                                                                       //                    enet_pll_outclk1.clk
		.enet_pll_outclk2_clk                            (),                                                                       //                    enet_pll_outclk2.clk
		.enet_pll_reset_reset                            (nios_cpu_qsys_inst_enet_pll_reset_bfm_reset_reset),                      //                      enet_pll_reset.reset
		.lcd_external_RS                                 (nios_cpu_qsys_inst_lcd_external_rs),                                     //                        lcd_external.RS
		.lcd_external_RW                                 (nios_cpu_qsys_inst_lcd_external_rw),                                     //                                    .RW
		.lcd_external_data                               (nios_cpu_qsys_inst_lcd_external_data),                                   //                                    .data
		.lcd_external_E                                  (nios_cpu_qsys_inst_lcd_external_e),                                      //                                    .E
		.merged_resets_in_reset_reset_n                  (nios_cpu_qsys_inst_merged_resets_in_reset_bfm_reset_reset),              //              merged_resets_in_reset.reset_n
		.samplenum_out_export                            (nios_cpu_qsys_inst_samplenum_out_export),                                //                       samplenum_out.export
		.tse_mac_mac_mdio_connection_mdc                 (nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdc),                     //         tse_mac_mac_mdio_connection.mdc
		.tse_mac_mac_mdio_connection_mdio_in             (nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_bfm_conduit_mdio_in),     //                                    .mdio_in
		.tse_mac_mac_mdio_connection_mdio_out            (nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdio_out),                //                                    .mdio_out
		.tse_mac_mac_mdio_connection_mdio_oen            (nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdio_oen),                //                                    .mdio_oen
		.tse_mac_mac_rgmii_connection_rgmii_in           (nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_bfm_conduit_rgmii_in),   //        tse_mac_mac_rgmii_connection.rgmii_in
		.tse_mac_mac_rgmii_connection_rgmii_out          (nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_rgmii_out),              //                                    .rgmii_out
		.tse_mac_mac_rgmii_connection_rx_control         (nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_bfm_conduit_rx_control), //                                    .rx_control
		.tse_mac_mac_rgmii_connection_tx_control         (nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_tx_control),             //                                    .tx_control
		.tse_mac_mac_status_connection_set_10            (nios_cpu_qsys_inst_tse_mac_mac_status_connection_bfm_conduit_set_10),    //       tse_mac_mac_status_connection.set_10
		.tse_mac_mac_status_connection_set_1000          (nios_cpu_qsys_inst_tse_mac_mac_status_connection_bfm_conduit_set_1000),  //                                    .set_1000
		.tse_mac_mac_status_connection_eth_mode          (nios_cpu_qsys_inst_tse_mac_mac_status_connection_eth_mode),              //                                    .eth_mode
		.tse_mac_mac_status_connection_ena_10            (nios_cpu_qsys_inst_tse_mac_mac_status_connection_ena_10),                //                                    .ena_10
		.tse_mac_pcs_mac_rx_clock_connection_clk         (nios_cpu_qsys_inst_tse_mac_pcs_mac_rx_clock_connection_bfm_clk_clk),     // tse_mac_pcs_mac_rx_clock_connection.clk
		.tse_mac_pcs_mac_tx_clock_connection_clk         (nios_cpu_qsys_inst_tse_mac_pcs_mac_tx_clock_connection_bfm_clk_clk),     // tse_mac_pcs_mac_tx_clock_connection.clk
		.wavesample_in_export                            (nios_cpu_qsys_inst_wavesample_in_bfm_conduit_export)                     //                       wavesample_in.export
	);

	altera_conduit_bfm nios_cpu_qsys_inst_adc_control_out_bfm (
		.sig_export (nios_cpu_qsys_inst_adc_control_out_export)  // conduit.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nios_cpu_qsys_inst_clk_bfm (
		.clk (nios_cpu_qsys_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm_0002 nios_cpu_qsys_inst_enet_pll_locked_bfm (
		.sig_export (nios_cpu_qsys_inst_enet_pll_locked_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (1),
		.INITIAL_RESET_CYCLES (50)
	) nios_cpu_qsys_inst_enet_pll_reset_bfm (
		.reset (nios_cpu_qsys_inst_enet_pll_reset_bfm_reset_reset), // reset.reset
		.clk   (nios_cpu_qsys_inst_clk_bfm_clk_clk)                 //   clk.clk
	);

	altera_conduit_bfm_0003 nios_cpu_qsys_inst_lcd_external_bfm (
		.sig_RS   (nios_cpu_qsys_inst_lcd_external_rs),   // conduit.RS
		.sig_RW   (nios_cpu_qsys_inst_lcd_external_rw),   //        .RW
		.sig_data (nios_cpu_qsys_inst_lcd_external_data), //        .data
		.sig_E    (nios_cpu_qsys_inst_lcd_external_e)     //        .E
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) nios_cpu_qsys_inst_merged_resets_in_reset_bfm (
		.reset (nios_cpu_qsys_inst_merged_resets_in_reset_bfm_reset_reset), // reset.reset_n
		.clk   (nios_cpu_qsys_inst_clk_bfm_clk_clk)                         //   clk.clk
	);

	altera_conduit_bfm_0004 nios_cpu_qsys_inst_samplenum_out_bfm (
		.sig_export (nios_cpu_qsys_inst_samplenum_out_export)  // conduit.export
	);

	altera_conduit_bfm_0005 nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_bfm (
		.sig_mdc      (nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdc),                 // conduit.mdc
		.sig_mdio_in  (nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_bfm_conduit_mdio_in), //        .mdio_in
		.sig_mdio_out (nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdio_out),            //        .mdio_out
		.sig_mdio_oen (nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdio_oen)             //        .mdio_oen
	);

	altera_conduit_bfm_0006 nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_bfm (
		.sig_rgmii_in   (nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_bfm_conduit_rgmii_in),   // conduit.rgmii_in
		.sig_rgmii_out  (nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_rgmii_out),              //        .rgmii_out
		.sig_rx_control (nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_bfm_conduit_rx_control), //        .rx_control
		.sig_tx_control (nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_tx_control)              //        .tx_control
	);

	altera_conduit_bfm_0007 nios_cpu_qsys_inst_tse_mac_mac_status_connection_bfm (
		.sig_set_10   (nios_cpu_qsys_inst_tse_mac_mac_status_connection_bfm_conduit_set_10),   // conduit.set_10
		.sig_set_1000 (nios_cpu_qsys_inst_tse_mac_mac_status_connection_bfm_conduit_set_1000), //        .set_1000
		.sig_eth_mode (nios_cpu_qsys_inst_tse_mac_mac_status_connection_eth_mode),             //        .eth_mode
		.sig_ena_10   (nios_cpu_qsys_inst_tse_mac_mac_status_connection_ena_10)                //        .ena_10
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nios_cpu_qsys_inst_tse_mac_pcs_mac_rx_clock_connection_bfm (
		.clk (nios_cpu_qsys_inst_tse_mac_pcs_mac_rx_clock_connection_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nios_cpu_qsys_inst_tse_mac_pcs_mac_tx_clock_connection_bfm (
		.clk (nios_cpu_qsys_inst_tse_mac_pcs_mac_tx_clock_connection_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm_0008 nios_cpu_qsys_inst_wavesample_in_bfm (
		.sig_export (nios_cpu_qsys_inst_wavesample_in_bfm_conduit_export)  // conduit.export
	);

	altera_tristate_conduit_bridge_translator cfi_flash_atb_bridge_0_tcb_translator (
		.in_tcm_address_out      (nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_address_out),      //  in.tcm_address_out
		.in_tcm_read_n_out       (nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_read_n_out),       //    .tcm_read_n_out
		.in_tcm_write_n_out      (nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_write_n_out),      //    .tcm_write_n_out
		.in_tcm_data_out         (nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_data_out),         //    .tcm_data_out
		.in_tcm_chipselect_n_out (nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out), //    .tcm_chipselect_n_out
		.tcm_address_out         (cfi_flash_atb_bridge_0_tcb_translator_out_tcm_address_out),          // out.tcm_address_out
		.tcm_read_n_out          (cfi_flash_atb_bridge_0_tcb_translator_out_tcm_read_n_out),           //    .tcm_read_n_out
		.tcm_write_n_out         (cfi_flash_atb_bridge_0_tcb_translator_out_tcm_write_n_out),          //    .tcm_write_n_out
		.tcm_data_out            (cfi_flash_atb_bridge_0_tcb_translator_out_tcm_data_out),             //    .tcm_data_out
		.tcm_chipselect_n_out    (cfi_flash_atb_bridge_0_tcb_translator_out_tcm_chipselect_n_out)      //    .tcm_chipselect_n_out
	);

	altera_conduit_bfm_0009 cfi_flash_atb_bridge_0_tcb_translator_out_bfm (
		.sig_tcm_address_out      (cfi_flash_atb_bridge_0_tcb_translator_out_tcm_address_out),      // conduit.tcm_address_out
		.sig_tcm_read_n_out       (cfi_flash_atb_bridge_0_tcb_translator_out_tcm_read_n_out),       //        .tcm_read_n_out
		.sig_tcm_write_n_out      (cfi_flash_atb_bridge_0_tcb_translator_out_tcm_write_n_out),      //        .tcm_write_n_out
		.sig_tcm_data_out         (cfi_flash_atb_bridge_0_tcb_translator_out_tcm_data_out),         //        .tcm_data_out
		.sig_tcm_chipselect_n_out (cfi_flash_atb_bridge_0_tcb_translator_out_tcm_chipselect_n_out)  //        .tcm_chipselect_n_out
	);

endmodule
