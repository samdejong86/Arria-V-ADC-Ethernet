// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
GMoGrLvGhUHYI1Rv5W0mjn6pCmKkAIWnmxmUAi7LNnRNiBxQHJldDbx7lmBP31lj
8TiRdQNandBUzCRn+TR5Hp88yvsB0wI13mmPQuFWHF/HajIxZR15zlONiGe8i+Vb
MywPo0nQh80zNxknCxcElUJnF/ArM44vD1zjqnnMCtF4lWeYbvEjQA==
//pragma protect end_key_block
//pragma protect digest_block
Oi9aTaFGqMQlyRyeCa74xN34BFc=
//pragma protect end_digest_block
//pragma protect data_block
X2iiEsPm4dXRP1qqrtr3HH+X9JJawqPaE+/MKoyCpcb3OjfKSchJgaa4iwN/vdbP
OnrR2NCnrQWShuOLpwf/Plm29RALEMB6hFVJnoi9jHRv8uQF/r8Rt8mmE93VqPoY
hq/uGwxTd5dPVB/C6XaK0SXa8aWZJGZWeooiCvqCNkvsjp0BcVfA5nylHpDAjhuh
ltdxt4/syFEg71xWoR1EvxwaNT3pbaSZhRJEdLyKPLBslaqs9h/GIPkkLyUAao6I
6RjR9Uclz8fkKPt/ATxnmVlLGdrB61ih14IKpUWFYCxvimsNVkGp63wLR+M9V09N
Rb8aTBFQA6SerTQ6LHX8JuWvzoKByR+WjA1iTHrmMLXGJnQ0JI08gin1atZG3Qb9
6XdrOJ7NAucjx4YJWAL0eQIMu1xyyhWb5SOAaBEwbGTQTQPXKh0t2Er1MkmxFVQ/
JEgNdbxR7flaFaCsd5xUmuYsB1XevazJoGqfQqgaWaQPx+rcE1ov+gWJUL/Olm+n
tLqdPsw9tV4MKS9hXhbniO13/Mtt0+xVhgMmbZrNeA1IzOLUcNS7owflTclmsYld
2nm1aMTAK0KlgTqq5nUAMHIzXihdfRjOjrljOnHZTBHadhv05fq/lS75GElvnQi8
/cMmry0nyNtJLbboEGPmZxR3sGCbAOsVDIx/8WOHYLvZ/WS9a0K7VAmAXe7zYw1K
+Kh66gW4FGM+0xw2uJZ6/TcOohW/oDYyp37zSrUPifcNX7E3B7acyTUIbgfyh4SV
igg/kBdtDMj4dP7E52MpscesH6TnwrFBKVLIpR6nFQXJwe5FzGFexUivqyCsi3BE
3+StpfYWdnqb/AijjsHruxZAyxdwhV6ZrNGW0H0DyqnuTblWFxu8QXSimXHzy6KX
sbCzVnfg3ARROVOfJ1ZWYqQlsKpNzJyortZMo+JXEPS4BP67JYDLCw4XWY+95n82
ddigHcF2wzqpJsIXcLY/o1TAqFF4CdQyZJmyOySxEbPEyPB6y3w61Ww1hPErZV0k
cYxasJRotXBTlKkEBav1/GifT7qWlgAVraXRAp9zSEUOWk0oX8VIoFP4a7HTArwB
Ph15B7mNkhPJFNYw2f7u8Yu042ALxUfJlmkz7Z/tJUX835E9iknLe8Vma+0GA0/f
Fbxn6T9hkUfocQ8/SDPxQU44OkYRfjJWedvFPMAXIyFMsD2uXoCKZzTleYwQe6t7
4hF2Nrl3N2rDsz3ZWKwsVTK7HyZgkzYpT+y56u6pwx87rjrZUcHf1SHrfO0IjqPB
4J7bEkiKbtv/COG3SUgXkuLiVU/4OBXY8/5R39W/ZWzJoVDO7nfCU0+h1CKwo5ey
R2dZKSxg1RAOD6Q2Z9ephbWCftRr/2MpbK5AcpApImeGvTc2v78+Gkf4OjtaIJji
/eXa0mabRMoFKtrM15VslSJNxnoc7xSKAcXz5p4EhZFCKv8GVq2xK6tR1VGAG19/
/nqFH6pCjqLqEUteSOsLx1isgs1bZGOM2TTLFoHer9lEOu+Dp+QUVLzQOPLwNS54
bwAjnRNOEm0DSzjj5DVuJ5cD4IO8fA6uMZ2zEPkNvHg3E8LGvtHsHpCfqLiXlFBx
lBF7ZmVc8Ndt5VmeprKHFyuimyimR72ecI6friguH2wc6d+ROZTnV2dPgSQTjOJY
oL7dxvwcBc14rrVi3a/alEAKpdzUplT4k5axxYeI2Eh0dbMZy6kjJXOO0TOWHoyC
fbXYIwEKzjPNPDrGs5AKgXQF22HNwnOJWlE3GoRqGk9WtQTjEbKjQayQVBiCUJG0
ALAOogsy4X06dW0wG34uFmJjvyi6AIZlfvJmo78IBVTnNzyesk4aGBpIePhWsvm/
rmWV7ImY8b8xrc+1Kau6xWfBPsBK7Vq4QDtPwuPjOxlRsMBQHAtW2fpbZCFXtZae
FIfzYn4jBfeSMOra8uZ5V3siTJ9YeAROXLgoGNktLjavNLAI58lvBFOa9iL5n1ov
+66MNvxvfyOGIhKPJKTHtGb44sS6KzTsBJmnn6Yeh/nBUtiUmY0GYh8JZDp8c5BW
syHaPNA8z3cxKrByL2Utcd2vb4o+3yxHhp9CbziaXqjJWu5HqtRRoC0LvLk0rITd
2OfKWdkjjh0T1rxH8gzXRMAeac6YFtKu8909VlThHWjyLTvdmPnPQZSRZlDAJ6PI
ZjV2L3yMwGXlCRd/WtnHr8UuT0OfjCo46Iica+lW5hK4TB8DXpDdtMu0sLViX9M6
J0ODh18H6/318lsHdZZd56gFzes0XVWD6cV4J8CQid+2AP5c3LXKtr1AYVUBkuK9
bw/fteNBZIBfnykYk74qudAq9EHXDHp0Y9a/GXW5pmPdGT00jb6IgTBhgAx+w12t
RXOjs0nnCMvKhYQPwbqZezPEuzy8o5PYtIV3kOPA85cES2h/iI6X1mfmQgKL+k1+
+1f9oXhqZr//YoaCzrJBWB4PxjPcRcqUOopHGQ8M0a6h0C7Zz8xfh29LJdlvTezI
Tywy19ZYL5vrURqeuRWIX4+Pr9K67tlVxFbauFY0Y3J2CnTeT/4uDTbPp0sYvE82
mGGCVVeew0aHyujX2avFdvoEE1LQZ1oNs613LPrde44/GoAyzMLwj7zYpuO2KBqy
6u9bF/3OceZFlG7KW8BoHprNRFqXK1edz9ilWS3C3jlZBZFVejt1YLCd+wY/TYKm
U/WinY893tAsgoeJlB1EUHyrXFRxGqrkEKRlkW78+H7R+RTgbTgptYkgsd5Jo67b
prRyYsn2oL9K8/US+rN8RMoANx63XIyrAHy15VphqYuumLBvnhnwip1x0snEV5l+
ds/ozFNJSYoIWaVj2vtXaxiM4RYBB5XbkIZ/CBr+HWTAEtK9VXyfJ5TEOoC0ug3+
BdoThJs0uaGcghtQf3XQBHdmtFUF7PXCSq6nQW73/IRcBxzjJ8BenlA+HZE0Rd3J
9BPO3BJgk5+b9Imqs1MMny2//kbrE8r+yocyNJl/itt/w6xAgg5Zs2VJVAfPQggV
hl0nEpl+4JeZ7/A1buokwiJ6M05Um0vLhXRHjWjUYLih7trGWsHbX5frLMjVwAyb
6sBRCjU9e1yhsN9nzGB/9XteWZGc4VCIJRapWm3ShD2xhUJ/NwLFvKGEq0UrJszS
2JmGwyXY58yox4F6J7d8SU94HZ7lftI1F0n6pnvFR/asQsmW5MaX18Iomd0MVGqB
kKnzih2SBlcJ5uMPX6OOdmndvpYPxFTUsdZP70AXA/h8RxWJb3ruC+n+x8i7ytfW
ho2s7oVi3METkigNNFVASJJuqYvQq6Fdr0gXDHXdU+dqY69HoRlTkdTq/KCHy3mj
CcYLe7Xi7D6f+OLT1OX3lvLpyEr5rDQAQIWAUa/Y1PqKN6Lg761T9c0fK49RMJ1q
+Tcg2ID8CX1iJ0ZyyumWw9kw6dlbrlF3fulai6uy6yz+8wuY9pu1IYNMHSLjIttv
EKC3lBSSY83jzh8Cw6VItMAwuhqxtfnzOK+YfF8mAZqM5DQJ0sSN9h9BoDYjXrpz
M9sGlgUoOqRzZ3NJ/AoB7oMt9zKfbkIldZ73cqDUMKYcEa2Blhbqf1x6Y3gP/lJm
aLebVY5C2xsnwHbEiVBgWLLNISLlFbn+wdRxtr84qXKyHkpkIzCQMVCVKecuau24
PjzGeumlNAOj+NCIdpeiZqvWVDCf6AK8/YMWAOxRrGBYQjywZep0W4Q5sYPilw/V
eNKjt+3xaq9kTB17TEHDmXr2pVJj7pH+bE0PjlfaE2TI3eEOQavY8v4WhApBbgmd
Y2bFdoVYyeS09QyRXAT8y91PBlU9ZBKeGT3JyxTOHJlurmbuQuKJHTnsTioZp383
aD64MqJI9HaKW6PFq5DWwyTmM3hs3ko9s/fRp0W+x1d7RMz+SfqaAW2L0Uq3vqCx
iUe1ZdkoeZKQR72s8obbEvpVNhobIA8fQebs+0Vjhk++3HnsNCFPW6Or8tBhgk7s
iDn+nxu1oLg83z4sLB2xvsaXaQaJ0UoZ/VeWUsFJ1BlU31Fp5IFu8OYSJ9Xw6NAY
besVa8OvJLNtqWnrllprjCYoMVPD9vtgTEdAvQROlsq2SdiYeqdG/F89vREAWgfD
/htxRzVEXFhu7sKmGD/KeoMGotNOOuxcQO7NEzrI5IMye3UEoZ5/ZCD8MGw1P/gA
10Q+MAMtZh3FwegkKxznFRRBwlAEOqt35GERra89T6iaAoo7HHOxFWJIFBzjlHGy
HyyRAGOqg5pq50grqIkdnVkmBPhbXh71MPC1B30GOv/GEAGhc8jmWoNWwUBUvGa5
WZO8VupDMad/amnnKnVP955T2Gd8iBsOEhKIodzeBF/ME/JdW6ETmtyyFojYdefg
YFmsIu7VWjIe5Gds7g7LWWSI7y0TweN+WPPF2q16D/uJiFCx4tDUVrX/Omw96q0F
LP+82ZgZjva0mjg8NTzdAE5FVh4Jrw5qUeNRAcDqwoSVcbrI+dVKTNDCfEBOMVtl
s/BVnJyv9TFiUv6Gu2Qdh6yiAwxsMLEIAG/mcog7sL6+ZxPuvipeOklvlLHZsN+B
6YwHNzgjRX/spKl9lB3juSI8frnfZLRsK+u+m6Uaev68fvEDmodXS3OYe0aJWwvE
KqM40d3ix3okRAc20Q9iQaJ622DZ3ZPaKlB935djZ/RMfEBBnSD+QFbFOGKAU256
fex5yhlWuP9S4OSrsqnweX7xM/dTfIDrgeynIJPbkUH5AO4RlaBIYAbJ5ZcOf0n/
hhQYoiPq8CzrpeQU11IqqOEh1M40tksbfpwx6dX1BmBfweKGzmxHTeaF/surMKOr
LE1Nn3kS1dJtW97H0UruJTYqc+D0UUlYCj8V6j4RLGSq0hR8QTHkI+HjpkSs4SNX
Lqu+nssyEyvX43k4eGdkt8U1smBQOzmS23B7ubLavvgd/ec6Xi4OTfh/V1rKKGnm
tewIrZUrQU99aSodmgMBNtvNnIl+7JzoHltzEl3CRycA2LLwABD6vSuLfMAqqID3
fcJ1lh4dUlsYoyMzyYzGwq457K7ZKjzSO8Z700p8KXFlvZ0NO6siHs7N3z7tWxXl
8K3SGsjzna6LkEOot+VBcNbERmU5H3jQPpNsDdgr8ocD2jt3ctTrZik19w9xZf4u
oiMEM0TcixvqRil96GdDCC4ELNAzpv0K1u7jHbVWsplOI8JIcjuo8ugzLaUMP6OR
FL5W9y2PntuqN+gEBIXhLeuxCNubk5BPD7PGgY21Rl1jfGfIKNJ/IO6f8dUDV7fY
FtPy9rfR5agM6+Y1rTJxU/hpubNW4HMx3XOvTAKTH6FIkmE3UXrZ8Dj8LMxwp0R3
PGS0H3BVHuuYKGtXGy+sx0ZWnycx8FFkGni2SVkHR8LUUfu/Ayhuqiffls+2uBpN
QmpXqoWJKNmXZv4isy+QXQRAKt30urlnubi/aAAnJNrWCImWKlH+0JKTmJcfpsb8
Ncx86vyL5kOgclMAJOHer+u7a3OWN9kEOfFM+ib/j5BrqCHUevQoUn1rWSYRB2y5
u8yOcN4WnO6p+TPlqiZzR259nIWMRLlL0e16+4WedU+dqr09qsQjhfgF2fHR8kWj
4w5pw177aoZQkiS1zSGYKx6rVyAYzZAsLq6BbefqgZKX5wV5f80SUht14/VEVYfM
v92tDg3aeTXLoe3RJ69mjNkEZuW95kdaru/q7h8i+pbLkFnw6DqXy6juiz3CRsnC
hjaDjIuSNbZTuViQwmlv1YRaI554NEN+IZGAb/hdjZBdsbAjuGxmrC6jqwR2LLDP
isFAivexehItBEyUi4DsdvmHc16yAGzJUSa+E2oQ2Hs54LomshlY3S6bd4CIjz0h
ah4zoxaxXGpthlw5SOzDva8/omJtW0Z6jK5n9jB/AfLP119RhmukKyTPcXBwkM5R
+taEyPtnF44bh4RLRRDIJyoL8ZMsTVtSyDJTBlY/Xg5GMfL9pvQSUTsodxG2dMgc
5JQtAibck5M5G4zcomsGI2VL7pyP+WFd40N9rWdtXOy9Bw1CCfgeNyoNJqa2eDXU
LPaGJfZF2ijHzHQD44wD+daMzVRK+TVvOLP3TgKIwlUHAAbrWegQXtajFTMSGR3G
Qi7YzJmZ1yb2MlH28ZF+oeDcwUfFZ8QKkK+gR/6KXeim49kpvIIUK33nHbKpVM7B
InKA+OCscv0oatpkvHgKVBrQcG9tom+wiEAag6V/4kVSJs0+PF4NeXdEkXMvsDhF
yvJybAK/tsltB94/FCuT8cnpFv5ihwUDoVjHIAlMpBY7KgWnOOSbIqXFnTBETXoQ
rM58Ibyvyu3DKKriHR4qccu8iHFlfbe1dlIVp1QZgafUFhK9Y9+W1i1/BN9BKBeu
Id/b40CrQ1yhyTphAIT4tSPie4whpjsCh/pOfsABZG5eVlpmnpy46881dPDL0OMF
ydaQyOgm3RSS9LjfEmRtxvLqh/P6Z8n+uc5ANGbNEgiJdK9+/x9jzYejdbp8HVYj
SsqI4DSykt+erZnnJhXgM7Rlh/9PjvpQQoE/C7PCRMwqpYUtltJEmf4eeSAxBVQF
/gzglRNnLAcDKgIDm/mTVLU1LODnORk2zKHfjo9J1WS1QcaNlCGnl1NSv2P193ai
HmpkdmNXOEFYisZom4e/xflQ/svvfre+Peb3UDWLs5Ns9WnQ5KYkK8kzY2AjMFda
85V8r2gdwTF5PkJsK79dvT/sS8k94vkH07+KdFn7JRGEtEET4edMQaPlQDAcHU2O
RnsXNsSk6HmptFhM69i7KoXJRbM3nec+TwSNgWmuTVYEo1W4iIbs/Ex/znKwKL/m
g5JHY5UQUHBYJVkoGNmsVsQ0Wrz2XXpQNXF5ANmu0tlV1/dfrsLDmu5qVKVCbnjQ
pqcpw9hdFAuKgubbxIGxkQbK0b6XAvZRamQ8rwryzaJo4sa2F7O48ryJLaCy7try
NLZ7AU3ZPc5XeG0tiDD68ozDKFbbqg9tppOYm7FvhaNkJKyhVo849uVyp1nogW4W
KqpsHws0Z1JUOQ/3EmwlxYZoZ3hDUgeCj/OTGlnovQhCoxWy412IJJz2WoW6fChk
h6YQbMSoN6FKOiRsEy0SBjJ1MDsZyekRiH3912CTzq4xvNblxDZ8A2PqZcVJGoP0

//pragma protect end_data_block
//pragma protect digest_block
UfMYsF9+Ycks8qbwx8pZ/drMH1A=
//pragma protect end_digest_block
//pragma protect end_protected
