-- Nios_CPU_qsys_tb.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Nios_CPU_qsys_tb is
end entity Nios_CPU_qsys_tb;

architecture rtl of Nios_CPU_qsys_tb is
	component Nios_CPU_qsys is
		port (
			adc_control_out_export                          : out   std_logic_vector(7 downto 0);                     -- export
			cfi_flash_atb_bridge_0_out_tcm_address_out      : out   std_logic_vector(26 downto 0);                    -- tcm_address_out
			cfi_flash_atb_bridge_0_out_tcm_read_n_out       : out   std_logic_vector(0 downto 0);                     -- tcm_read_n_out
			cfi_flash_atb_bridge_0_out_tcm_write_n_out      : out   std_logic_vector(0 downto 0);                     -- tcm_write_n_out
			cfi_flash_atb_bridge_0_out_tcm_data_out         : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out : out   std_logic_vector(0 downto 0);                     -- tcm_chipselect_n_out
			clk_clk                                         : in    std_logic                     := 'X';             -- clk
			enet_pll_locked_export                          : out   std_logic;                                        -- export
			enet_pll_outclk0_clk                            : out   std_logic;                                        -- clk
			enet_pll_outclk1_clk                            : out   std_logic;                                        -- clk
			enet_pll_outclk2_clk                            : out   std_logic;                                        -- clk
			enet_pll_reset_reset                            : in    std_logic                     := 'X';             -- reset
			lcd_external_RS                                 : out   std_logic;                                        -- RS
			lcd_external_RW                                 : out   std_logic;                                        -- RW
			lcd_external_data                               : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			lcd_external_E                                  : out   std_logic;                                        -- E
			merged_resets_in_reset_reset_n                  : in    std_logic                     := 'X';             -- reset_n
			samplenum_out_export                            : out   std_logic_vector(15 downto 0);                    -- export
			tse_mac_mac_mdio_connection_mdc                 : out   std_logic;                                        -- mdc
			tse_mac_mac_mdio_connection_mdio_in             : in    std_logic                     := 'X';             -- mdio_in
			tse_mac_mac_mdio_connection_mdio_out            : out   std_logic;                                        -- mdio_out
			tse_mac_mac_mdio_connection_mdio_oen            : out   std_logic;                                        -- mdio_oen
			tse_mac_mac_rgmii_connection_rgmii_in           : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- rgmii_in
			tse_mac_mac_rgmii_connection_rgmii_out          : out   std_logic_vector(3 downto 0);                     -- rgmii_out
			tse_mac_mac_rgmii_connection_rx_control         : in    std_logic                     := 'X';             -- rx_control
			tse_mac_mac_rgmii_connection_tx_control         : out   std_logic;                                        -- tx_control
			tse_mac_mac_status_connection_set_10            : in    std_logic                     := 'X';             -- set_10
			tse_mac_mac_status_connection_set_1000          : in    std_logic                     := 'X';             -- set_1000
			tse_mac_mac_status_connection_eth_mode          : out   std_logic;                                        -- eth_mode
			tse_mac_mac_status_connection_ena_10            : out   std_logic;                                        -- ena_10
			tse_mac_pcs_mac_rx_clock_connection_clk         : in    std_logic                     := 'X';             -- clk
			tse_mac_pcs_mac_tx_clock_connection_clk         : in    std_logic                     := 'X';             -- clk
			wavesample_in_export                            : in    std_logic_vector(15 downto 0) := (others => 'X')  -- export
		);
	end component Nios_CPU_qsys;

	component altera_conduit_bfm is
		port (
			sig_export : in std_logic_vector(7 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_conduit_bfm_0002 is
		port (
			sig_export : in std_logic_vector(0 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0002;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_conduit_bfm_0003 is
		port (
			sig_RS   : in    std_logic_vector(0 downto 0) := (others => 'X'); -- RS
			sig_RW   : in    std_logic_vector(0 downto 0) := (others => 'X'); -- RW
			sig_data : inout std_logic_vector(7 downto 0) := (others => 'X'); -- data
			sig_E    : in    std_logic_vector(0 downto 0) := (others => 'X')  -- E
		);
	end component altera_conduit_bfm_0003;

	component altera_conduit_bfm_0004 is
		port (
			sig_export : in std_logic_vector(15 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0004;

	component altera_conduit_bfm_0005 is
		port (
			sig_mdc      : in  std_logic_vector(0 downto 0) := (others => 'X'); -- mdc
			sig_mdio_in  : out std_logic_vector(0 downto 0);                    -- mdio_in
			sig_mdio_out : in  std_logic_vector(0 downto 0) := (others => 'X'); -- mdio_out
			sig_mdio_oen : in  std_logic_vector(0 downto 0) := (others => 'X')  -- mdio_oen
		);
	end component altera_conduit_bfm_0005;

	component altera_conduit_bfm_0006 is
		port (
			sig_rgmii_in   : out std_logic_vector(3 downto 0);                    -- rgmii_in
			sig_rgmii_out  : in  std_logic_vector(3 downto 0) := (others => 'X'); -- rgmii_out
			sig_rx_control : out std_logic_vector(0 downto 0);                    -- rx_control
			sig_tx_control : in  std_logic_vector(0 downto 0) := (others => 'X')  -- tx_control
		);
	end component altera_conduit_bfm_0006;

	component altera_conduit_bfm_0007 is
		port (
			sig_set_10   : out std_logic_vector(0 downto 0);                    -- set_10
			sig_set_1000 : out std_logic_vector(0 downto 0);                    -- set_1000
			sig_eth_mode : in  std_logic_vector(0 downto 0) := (others => 'X'); -- eth_mode
			sig_ena_10   : in  std_logic_vector(0 downto 0) := (others => 'X')  -- ena_10
		);
	end component altera_conduit_bfm_0007;

	component altera_conduit_bfm_0008 is
		port (
			sig_export : out std_logic_vector(15 downto 0)   -- export
		);
	end component altera_conduit_bfm_0008;

	component altera_tristate_conduit_bridge_translator is
		port (
			in_tcm_address_out      : in    std_logic_vector(26 downto 0) := (others => 'X'); -- tcm_address_out
			in_tcm_read_n_out       : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tcm_read_n_out
			in_tcm_write_n_out      : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tcm_write_n_out
			in_tcm_data_out         : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			in_tcm_chipselect_n_out : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tcm_chipselect_n_out
			tcm_address_out         : out   std_logic_vector(26 downto 0);                    -- tcm_address_out
			tcm_read_n_out          : out   std_logic_vector(0 downto 0);                     -- tcm_read_n_out
			tcm_write_n_out         : out   std_logic_vector(0 downto 0);                     -- tcm_write_n_out
			tcm_data_out            : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			tcm_chipselect_n_out    : out   std_logic_vector(0 downto 0)                      -- tcm_chipselect_n_out
		);
	end component altera_tristate_conduit_bridge_translator;

	component altera_conduit_bfm_0009 is
		port (
			sig_tcm_address_out      : in    std_logic_vector(26 downto 0) := (others => 'X'); -- tcm_address_out
			sig_tcm_read_n_out       : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tcm_read_n_out
			sig_tcm_write_n_out      : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tcm_write_n_out
			sig_tcm_data_out         : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			sig_tcm_chipselect_n_out : in    std_logic_vector(0 downto 0)  := (others => 'X')  -- tcm_chipselect_n_out
		);
	end component altera_conduit_bfm_0009;

	signal nios_cpu_qsys_inst_clk_bfm_clk_clk                                     : std_logic;                     -- Nios_CPU_qsys_inst_clk_bfm:clk -> [Nios_CPU_qsys_inst:clk_clk, Nios_CPU_qsys_inst_enet_pll_reset_bfm:clk, Nios_CPU_qsys_inst_merged_resets_in_reset_bfm:clk]
	signal nios_cpu_qsys_inst_tse_mac_pcs_mac_rx_clock_connection_bfm_clk_clk     : std_logic;                     -- Nios_CPU_qsys_inst_tse_mac_pcs_mac_rx_clock_connection_bfm:clk -> Nios_CPU_qsys_inst:tse_mac_pcs_mac_rx_clock_connection_clk
	signal nios_cpu_qsys_inst_tse_mac_pcs_mac_tx_clock_connection_bfm_clk_clk     : std_logic;                     -- Nios_CPU_qsys_inst_tse_mac_pcs_mac_tx_clock_connection_bfm:clk -> Nios_CPU_qsys_inst:tse_mac_pcs_mac_tx_clock_connection_clk
	signal nios_cpu_qsys_inst_adc_control_out_export                              : std_logic_vector(7 downto 0);  -- Nios_CPU_qsys_inst:adc_control_out_export -> Nios_CPU_qsys_inst_adc_control_out_bfm:sig_export
	signal nios_cpu_qsys_inst_enet_pll_locked_export                              : std_logic;                     -- Nios_CPU_qsys_inst:enet_pll_locked_export -> Nios_CPU_qsys_inst_enet_pll_locked_bfm:sig_export
	signal nios_cpu_qsys_inst_lcd_external_rs                                     : std_logic;                     -- Nios_CPU_qsys_inst:lcd_external_RS -> Nios_CPU_qsys_inst_lcd_external_bfm:sig_RS
	signal nios_cpu_qsys_inst_lcd_external_data                                   : std_logic_vector(7 downto 0);  -- [] -> [Nios_CPU_qsys_inst:lcd_external_data, Nios_CPU_qsys_inst_lcd_external_bfm:sig_data]
	signal nios_cpu_qsys_inst_lcd_external_rw                                     : std_logic;                     -- Nios_CPU_qsys_inst:lcd_external_RW -> Nios_CPU_qsys_inst_lcd_external_bfm:sig_RW
	signal nios_cpu_qsys_inst_lcd_external_e                                      : std_logic;                     -- Nios_CPU_qsys_inst:lcd_external_E -> Nios_CPU_qsys_inst_lcd_external_bfm:sig_E
	signal cfi_flash_atb_bridge_0_tcb_translator_out_tcm_chipselect_n_out         : std_logic_vector(0 downto 0);  -- cfi_flash_atb_bridge_0_tcb_translator:tcm_chipselect_n_out -> cfi_flash_atb_bridge_0_tcb_translator_out_bfm:sig_tcm_chipselect_n_out
	signal cfi_flash_atb_bridge_0_tcb_translator_out_tcm_address_out              : std_logic_vector(26 downto 0); -- cfi_flash_atb_bridge_0_tcb_translator:tcm_address_out -> cfi_flash_atb_bridge_0_tcb_translator_out_bfm:sig_tcm_address_out
	signal cfi_flash_atb_bridge_0_tcb_translator_out_tcm_data_out                 : std_logic_vector(15 downto 0); -- [] -> [cfi_flash_atb_bridge_0_tcb_translator:tcm_data_out, cfi_flash_atb_bridge_0_tcb_translator_out_bfm:sig_tcm_data_out]
	signal cfi_flash_atb_bridge_0_tcb_translator_out_tcm_read_n_out               : std_logic_vector(0 downto 0);  -- cfi_flash_atb_bridge_0_tcb_translator:tcm_read_n_out -> cfi_flash_atb_bridge_0_tcb_translator_out_bfm:sig_tcm_read_n_out
	signal cfi_flash_atb_bridge_0_tcb_translator_out_tcm_write_n_out              : std_logic_vector(0 downto 0);  -- cfi_flash_atb_bridge_0_tcb_translator:tcm_write_n_out -> cfi_flash_atb_bridge_0_tcb_translator_out_bfm:sig_tcm_write_n_out
	signal nios_cpu_qsys_inst_samplenum_out_export                                : std_logic_vector(15 downto 0); -- Nios_CPU_qsys_inst:samplenum_out_export -> Nios_CPU_qsys_inst_samplenum_out_bfm:sig_export
	signal nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_bfm_conduit_mdio_in     : std_logic_vector(0 downto 0);  -- Nios_CPU_qsys_inst_tse_mac_mac_mdio_connection_bfm:sig_mdio_in -> Nios_CPU_qsys_inst:tse_mac_mac_mdio_connection_mdio_in
	signal nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdio_oen                : std_logic;                     -- Nios_CPU_qsys_inst:tse_mac_mac_mdio_connection_mdio_oen -> Nios_CPU_qsys_inst_tse_mac_mac_mdio_connection_bfm:sig_mdio_oen
	signal nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdio_out                : std_logic;                     -- Nios_CPU_qsys_inst:tse_mac_mac_mdio_connection_mdio_out -> Nios_CPU_qsys_inst_tse_mac_mac_mdio_connection_bfm:sig_mdio_out
	signal nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdc                     : std_logic;                     -- Nios_CPU_qsys_inst:tse_mac_mac_mdio_connection_mdc -> Nios_CPU_qsys_inst_tse_mac_mac_mdio_connection_bfm:sig_mdc
	signal nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_tx_control             : std_logic;                     -- Nios_CPU_qsys_inst:tse_mac_mac_rgmii_connection_tx_control -> Nios_CPU_qsys_inst_tse_mac_mac_rgmii_connection_bfm:sig_tx_control
	signal nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_bfm_conduit_rx_control : std_logic_vector(0 downto 0);  -- Nios_CPU_qsys_inst_tse_mac_mac_rgmii_connection_bfm:sig_rx_control -> Nios_CPU_qsys_inst:tse_mac_mac_rgmii_connection_rx_control
	signal nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_bfm_conduit_rgmii_in   : std_logic_vector(3 downto 0);  -- Nios_CPU_qsys_inst_tse_mac_mac_rgmii_connection_bfm:sig_rgmii_in -> Nios_CPU_qsys_inst:tse_mac_mac_rgmii_connection_rgmii_in
	signal nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_rgmii_out              : std_logic_vector(3 downto 0);  -- Nios_CPU_qsys_inst:tse_mac_mac_rgmii_connection_rgmii_out -> Nios_CPU_qsys_inst_tse_mac_mac_rgmii_connection_bfm:sig_rgmii_out
	signal nios_cpu_qsys_inst_tse_mac_mac_status_connection_ena_10                : std_logic;                     -- Nios_CPU_qsys_inst:tse_mac_mac_status_connection_ena_10 -> Nios_CPU_qsys_inst_tse_mac_mac_status_connection_bfm:sig_ena_10
	signal nios_cpu_qsys_inst_tse_mac_mac_status_connection_eth_mode              : std_logic;                     -- Nios_CPU_qsys_inst:tse_mac_mac_status_connection_eth_mode -> Nios_CPU_qsys_inst_tse_mac_mac_status_connection_bfm:sig_eth_mode
	signal nios_cpu_qsys_inst_tse_mac_mac_status_connection_bfm_conduit_set_1000  : std_logic_vector(0 downto 0);  -- Nios_CPU_qsys_inst_tse_mac_mac_status_connection_bfm:sig_set_1000 -> Nios_CPU_qsys_inst:tse_mac_mac_status_connection_set_1000
	signal nios_cpu_qsys_inst_tse_mac_mac_status_connection_bfm_conduit_set_10    : std_logic_vector(0 downto 0);  -- Nios_CPU_qsys_inst_tse_mac_mac_status_connection_bfm:sig_set_10 -> Nios_CPU_qsys_inst:tse_mac_mac_status_connection_set_10
	signal nios_cpu_qsys_inst_wavesample_in_bfm_conduit_export                    : std_logic_vector(15 downto 0); -- Nios_CPU_qsys_inst_wavesample_in_bfm:sig_export -> Nios_CPU_qsys_inst:wavesample_in_export
	signal nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out     : std_logic_vector(0 downto 0);  -- Nios_CPU_qsys_inst:cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out -> cfi_flash_atb_bridge_0_tcb_translator:in_tcm_chipselect_n_out
	signal nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_address_out          : std_logic_vector(26 downto 0); -- Nios_CPU_qsys_inst:cfi_flash_atb_bridge_0_out_tcm_address_out -> cfi_flash_atb_bridge_0_tcb_translator:in_tcm_address_out
	signal nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_data_out             : std_logic_vector(15 downto 0); -- [] -> [Nios_CPU_qsys_inst:cfi_flash_atb_bridge_0_out_tcm_data_out, cfi_flash_atb_bridge_0_tcb_translator:in_tcm_data_out]
	signal nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_read_n_out           : std_logic_vector(0 downto 0);  -- Nios_CPU_qsys_inst:cfi_flash_atb_bridge_0_out_tcm_read_n_out -> cfi_flash_atb_bridge_0_tcb_translator:in_tcm_read_n_out
	signal nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_write_n_out          : std_logic_vector(0 downto 0);  -- Nios_CPU_qsys_inst:cfi_flash_atb_bridge_0_out_tcm_write_n_out -> cfi_flash_atb_bridge_0_tcb_translator:in_tcm_write_n_out
	signal nios_cpu_qsys_inst_enet_pll_reset_bfm_reset_reset                      : std_logic;                     -- Nios_CPU_qsys_inst_enet_pll_reset_bfm:reset -> Nios_CPU_qsys_inst:enet_pll_reset_reset
	signal nios_cpu_qsys_inst_merged_resets_in_reset_bfm_reset_reset              : std_logic;                     -- Nios_CPU_qsys_inst_merged_resets_in_reset_bfm:reset -> Nios_CPU_qsys_inst:merged_resets_in_reset_reset_n

begin

	nios_cpu_qsys_inst : component Nios_CPU_qsys
		port map (
			adc_control_out_export                          => nios_cpu_qsys_inst_adc_control_out_export,                                 --                     adc_control_out.export
			cfi_flash_atb_bridge_0_out_tcm_address_out      => nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_address_out,             --          cfi_flash_atb_bridge_0_out.tcm_address_out
			cfi_flash_atb_bridge_0_out_tcm_read_n_out       => nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_read_n_out,              --                                    .tcm_read_n_out
			cfi_flash_atb_bridge_0_out_tcm_write_n_out      => nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_write_n_out,             --                                    .tcm_write_n_out
			cfi_flash_atb_bridge_0_out_tcm_data_out         => nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_data_out,                --                                    .tcm_data_out
			cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out => nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out,        --                                    .tcm_chipselect_n_out
			clk_clk                                         => nios_cpu_qsys_inst_clk_bfm_clk_clk,                                        --                                 clk.clk
			enet_pll_locked_export                          => nios_cpu_qsys_inst_enet_pll_locked_export,                                 --                     enet_pll_locked.export
			enet_pll_outclk0_clk                            => open,                                                                      --                    enet_pll_outclk0.clk
			enet_pll_outclk1_clk                            => open,                                                                      --                    enet_pll_outclk1.clk
			enet_pll_outclk2_clk                            => open,                                                                      --                    enet_pll_outclk2.clk
			enet_pll_reset_reset                            => nios_cpu_qsys_inst_enet_pll_reset_bfm_reset_reset,                         --                      enet_pll_reset.reset
			lcd_external_RS                                 => nios_cpu_qsys_inst_lcd_external_rs,                                        --                        lcd_external.RS
			lcd_external_RW                                 => nios_cpu_qsys_inst_lcd_external_rw,                                        --                                    .RW
			lcd_external_data                               => nios_cpu_qsys_inst_lcd_external_data,                                      --                                    .data
			lcd_external_E                                  => nios_cpu_qsys_inst_lcd_external_e,                                         --                                    .E
			merged_resets_in_reset_reset_n                  => nios_cpu_qsys_inst_merged_resets_in_reset_bfm_reset_reset,                 --              merged_resets_in_reset.reset_n
			samplenum_out_export                            => nios_cpu_qsys_inst_samplenum_out_export,                                   --                       samplenum_out.export
			tse_mac_mac_mdio_connection_mdc                 => nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdc,                        --         tse_mac_mac_mdio_connection.mdc
			tse_mac_mac_mdio_connection_mdio_in             => nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_bfm_conduit_mdio_in(0),     --                                    .mdio_in
			tse_mac_mac_mdio_connection_mdio_out            => nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdio_out,                   --                                    .mdio_out
			tse_mac_mac_mdio_connection_mdio_oen            => nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdio_oen,                   --                                    .mdio_oen
			tse_mac_mac_rgmii_connection_rgmii_in           => nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_bfm_conduit_rgmii_in,      --        tse_mac_mac_rgmii_connection.rgmii_in
			tse_mac_mac_rgmii_connection_rgmii_out          => nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_rgmii_out,                 --                                    .rgmii_out
			tse_mac_mac_rgmii_connection_rx_control         => nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_bfm_conduit_rx_control(0), --                                    .rx_control
			tse_mac_mac_rgmii_connection_tx_control         => nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_tx_control,                --                                    .tx_control
			tse_mac_mac_status_connection_set_10            => nios_cpu_qsys_inst_tse_mac_mac_status_connection_bfm_conduit_set_10(0),    --       tse_mac_mac_status_connection.set_10
			tse_mac_mac_status_connection_set_1000          => nios_cpu_qsys_inst_tse_mac_mac_status_connection_bfm_conduit_set_1000(0),  --                                    .set_1000
			tse_mac_mac_status_connection_eth_mode          => nios_cpu_qsys_inst_tse_mac_mac_status_connection_eth_mode,                 --                                    .eth_mode
			tse_mac_mac_status_connection_ena_10            => nios_cpu_qsys_inst_tse_mac_mac_status_connection_ena_10,                   --                                    .ena_10
			tse_mac_pcs_mac_rx_clock_connection_clk         => nios_cpu_qsys_inst_tse_mac_pcs_mac_rx_clock_connection_bfm_clk_clk,        -- tse_mac_pcs_mac_rx_clock_connection.clk
			tse_mac_pcs_mac_tx_clock_connection_clk         => nios_cpu_qsys_inst_tse_mac_pcs_mac_tx_clock_connection_bfm_clk_clk,        -- tse_mac_pcs_mac_tx_clock_connection.clk
			wavesample_in_export                            => nios_cpu_qsys_inst_wavesample_in_bfm_conduit_export                        --                       wavesample_in.export
		);

	nios_cpu_qsys_inst_adc_control_out_bfm : component altera_conduit_bfm
		port map (
			sig_export => nios_cpu_qsys_inst_adc_control_out_export  -- conduit.export
		);

	nios_cpu_qsys_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => nios_cpu_qsys_inst_clk_bfm_clk_clk  -- clk.clk
		);

	nios_cpu_qsys_inst_enet_pll_locked_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export(0) => nios_cpu_qsys_inst_enet_pll_locked_export  -- conduit.export
		);

	nios_cpu_qsys_inst_enet_pll_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 1,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => nios_cpu_qsys_inst_enet_pll_reset_bfm_reset_reset, -- reset.reset
			clk   => nios_cpu_qsys_inst_clk_bfm_clk_clk                 --   clk.clk
		);

	nios_cpu_qsys_inst_lcd_external_bfm : component altera_conduit_bfm_0003
		port map (
			sig_RS(0) => nios_cpu_qsys_inst_lcd_external_rs,   -- conduit.RS
			sig_RW(0) => nios_cpu_qsys_inst_lcd_external_rw,   --        .RW
			sig_data  => nios_cpu_qsys_inst_lcd_external_data, --        .data
			sig_E(0)  => nios_cpu_qsys_inst_lcd_external_e     --        .E
		);

	nios_cpu_qsys_inst_merged_resets_in_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => nios_cpu_qsys_inst_merged_resets_in_reset_bfm_reset_reset, -- reset.reset_n
			clk   => nios_cpu_qsys_inst_clk_bfm_clk_clk                         --   clk.clk
		);

	nios_cpu_qsys_inst_samplenum_out_bfm : component altera_conduit_bfm_0004
		port map (
			sig_export => nios_cpu_qsys_inst_samplenum_out_export  -- conduit.export
		);

	nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_bfm : component altera_conduit_bfm_0005
		port map (
			sig_mdc(0)      => nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdc,                 -- conduit.mdc
			sig_mdio_in     => nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_bfm_conduit_mdio_in, --        .mdio_in
			sig_mdio_out(0) => nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdio_out,            --        .mdio_out
			sig_mdio_oen(0) => nios_cpu_qsys_inst_tse_mac_mac_mdio_connection_mdio_oen             --        .mdio_oen
		);

	nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_bfm : component altera_conduit_bfm_0006
		port map (
			sig_rgmii_in      => nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_bfm_conduit_rgmii_in,   -- conduit.rgmii_in
			sig_rgmii_out     => nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_rgmii_out,              --        .rgmii_out
			sig_rx_control    => nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_bfm_conduit_rx_control, --        .rx_control
			sig_tx_control(0) => nios_cpu_qsys_inst_tse_mac_mac_rgmii_connection_tx_control              --        .tx_control
		);

	nios_cpu_qsys_inst_tse_mac_mac_status_connection_bfm : component altera_conduit_bfm_0007
		port map (
			sig_set_10      => nios_cpu_qsys_inst_tse_mac_mac_status_connection_bfm_conduit_set_10,   -- conduit.set_10
			sig_set_1000    => nios_cpu_qsys_inst_tse_mac_mac_status_connection_bfm_conduit_set_1000, --        .set_1000
			sig_eth_mode(0) => nios_cpu_qsys_inst_tse_mac_mac_status_connection_eth_mode,             --        .eth_mode
			sig_ena_10(0)   => nios_cpu_qsys_inst_tse_mac_mac_status_connection_ena_10                --        .ena_10
		);

	nios_cpu_qsys_inst_tse_mac_pcs_mac_rx_clock_connection_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => nios_cpu_qsys_inst_tse_mac_pcs_mac_rx_clock_connection_bfm_clk_clk  -- clk.clk
		);

	nios_cpu_qsys_inst_tse_mac_pcs_mac_tx_clock_connection_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => nios_cpu_qsys_inst_tse_mac_pcs_mac_tx_clock_connection_bfm_clk_clk  -- clk.clk
		);

	nios_cpu_qsys_inst_wavesample_in_bfm : component altera_conduit_bfm_0008
		port map (
			sig_export => nios_cpu_qsys_inst_wavesample_in_bfm_conduit_export  -- conduit.export
		);

	cfi_flash_atb_bridge_0_tcb_translator : component altera_tristate_conduit_bridge_translator
		port map (
			in_tcm_address_out      => nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_address_out,      --  in.tcm_address_out
			in_tcm_read_n_out       => nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_read_n_out,       --    .tcm_read_n_out
			in_tcm_write_n_out      => nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_write_n_out,      --    .tcm_write_n_out
			in_tcm_data_out         => nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_data_out,         --    .tcm_data_out
			in_tcm_chipselect_n_out => nios_cpu_qsys_inst_cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out, --    .tcm_chipselect_n_out
			tcm_address_out         => cfi_flash_atb_bridge_0_tcb_translator_out_tcm_address_out,          -- out.tcm_address_out
			tcm_read_n_out          => cfi_flash_atb_bridge_0_tcb_translator_out_tcm_read_n_out,           --    .tcm_read_n_out
			tcm_write_n_out         => cfi_flash_atb_bridge_0_tcb_translator_out_tcm_write_n_out,          --    .tcm_write_n_out
			tcm_data_out            => cfi_flash_atb_bridge_0_tcb_translator_out_tcm_data_out,             --    .tcm_data_out
			tcm_chipselect_n_out    => cfi_flash_atb_bridge_0_tcb_translator_out_tcm_chipselect_n_out      --    .tcm_chipselect_n_out
		);

	cfi_flash_atb_bridge_0_tcb_translator_out_bfm : component altera_conduit_bfm_0009
		port map (
			sig_tcm_address_out      => cfi_flash_atb_bridge_0_tcb_translator_out_tcm_address_out,      -- conduit.tcm_address_out
			sig_tcm_read_n_out       => cfi_flash_atb_bridge_0_tcb_translator_out_tcm_read_n_out,       --        .tcm_read_n_out
			sig_tcm_write_n_out      => cfi_flash_atb_bridge_0_tcb_translator_out_tcm_write_n_out,      --        .tcm_write_n_out
			sig_tcm_data_out         => cfi_flash_atb_bridge_0_tcb_translator_out_tcm_data_out,         --        .tcm_data_out
			sig_tcm_chipselect_n_out => cfi_flash_atb_bridge_0_tcb_translator_out_tcm_chipselect_n_out  --        .tcm_chipselect_n_out
		);

end architecture rtl; -- of Nios_CPU_qsys_tb
