
module delayVec_vhdl(
	input [13:0] ADC_IN,
	input clk,
	output [13:0] DelayVec [100]
);
endmodule 